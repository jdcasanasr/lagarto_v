`define		riscv_pkg_XLEN						64
`define		change_pc							1:0
`define		instruction_memory_valid			43
`define		instruccion_memory_virtual_addres	42:3
`define		invalidate_icache					2
`define		invalidate_buffer					1
`define		invalidate_fecth					0
`define		fetch_o_pc							291:228
`define		fetch_o_resp_icache_cpu_i			227:196
`define		fetch_o_valid						195
`define		fetch_o_is_branch					194
`define		fetch_o_branch_decision				193
`define		fetch_o_branch_address				192-:`riscv_pkg_XLEN
`define		fetch_o_exception_cause				128:65
`define		fetch_o_exception_origin			64:1
`define		fetch_o_exception_valid				0
`define		branch_predictor_i_pc				129:66
`define		branch_predictor_i_adrres_result	65:2
`define		branch_predictor_i_taken_result		1
`define		branch_predictor_i_execution		0
`define		INSTR_ADDR_MISALIGNED				64'h0
`define		INSTR_ACCESS_FAULT					64'h1
`define		INSTR_PAGE_FAULT					64'hc