`define		instruction_length
`define		immediate_length
`define		
`define		
`define		
`define		
`define		
`define		
`define		
`define		
`define		
`define		