`define		not_request				2'b01
`define		request_valid			2'b10
`define		response_icache_data	32:1