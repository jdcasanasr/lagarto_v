`include	"Headers/riscv_vector.vh"
module shift_right(
	input			[2:0]		vsew_i,
	input			[127:0]	a,
	input			[127:0]	b,
	output reg	[127:0]	s
);
	
	always @(*)
		begin
			case(vsew_i)
				`vsew_8:
					begin
						s[7:0] 		<=	a[7:0]		>>		b[2:0];
						s[15:8]		<=	a[15:8]		>>		b[10:8];
						s[23:16]		<=	a[23:16]		>>		b[18:16];
						s[31:24]		<=	a[31:24]		>>		b[26:24];
						s[39:32]		<=	a[39:32]		>>		b[34:32];
						s[47:40]		<=	a[47:40]		>>		b[42:40];
						s[55:48]		<=	a[55:48]		>>		b[50:48];
						s[63:56]		<=	a[63:56]		>>		b[58:56];
						s[71:64]		<=	a[71:64]		>>		b[66:64];
						s[79:72]		<=	a[79:72]		>>		b[74:72];
						s[87:80]		<=	a[87:80]		>>		b[82:80];
						s[95:88]		<=	a[95:88]		>>		b[90:88];
						s[103:96]	<=	a[103:96]	>>		b[98:96];
						s[111:104]	<=	a[111:104]	>>		b[106:104];
						s[119:112]	<=	a[119:112]	>>		b[114:112];
						s[127:120]	<=	a[127:120]	>>		b[122:120];
					end
				`vsew_16:
					begin
						s[15:0] 		<=	a[15:0]		>>		b[3:0];
						s[31:16]		<=	a[31:16]		>>		b[19:16];
						s[47:32]		<=	a[47:32]		>>		b[35:32];
						s[63:48]		<=	a[63:48]		>>		b[51:48];
						s[79:64]		<=	a[79:64]		>>		b[67:64];
						s[95:80]		<=	a[95:80]		>>		b[83:80];
						s[111:96]	<=	a[111:96]	>>		b[99:96];
						s[127:112]	<=	a[127:112]	>>		b[115:112];
					end
				`vsew_32:
					begin
						s[31:0] 		<=	a[31:0] 		>>		b[4:0];
						s[63:32]		<=	a[63:32]		>>		b[36:32];
						s[95:64]		<=	a[95:64]		>>		b[68:64];
						s[127:96]	<=	a[127:96]	>>		b[100:96];
					end
				`vsew_64:
					begin
						s[63:0] 		<=	a[63:0] 		>>		b[5:0];
						s[127:64]	<=	a[127:64]	>>		b[69:64];
					end
				default:
						s <= 'b0;
			endcase
		end
endmodule 