`define lui_type 		7'b0110111
`define auipc_type 		7'b0010111
`define jal_type 		7'b1101111
`define jalr_type 		7'b1100111
`define branch_type 	7'b1100011
`define load_type 		7'b0000011
`define store_type 		7'b0100011
`define atomic_type 	7'b0101111
`define alu_i_type 		7'b0010011
`define alu_type 		7'b0110011
`define alu_i_w_type 	7'b0011011
`define alu_w_type 		7'b0111011
`define fence_type 		7'b0001111
`define system_type		7'b1110011		
