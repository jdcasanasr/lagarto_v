// Test Cases for the Vector Register File
// Read Vectors
`define read_vv
`define read_vx
`define read_vi

`define read_vv_vmask
`define read_vx_vmask
`define read_vi_vmask