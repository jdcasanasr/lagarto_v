// Reference: https://github.com/jdcasanasr/lagarto_v/tree/main/doc

/*	Resource Vectors
		System Vector
			BIT 5 	-> 	Cache Sync Atomic Operation (AMO)
			BIT 4 	-> 	System Operation (SYS)
			BIT 3 	-> 	Halt Operation (HALT)
			BIT 2 	-> 	Memory Sync Fence Operation (FENCE)
			BIT 1 	-> 	Memory Load Operation (L)
			BIT 0 	-> 	Memory Store Operation (S)
			
		Resource Vector
			BIT 21 	-> 	Vector Conversion Unit (VFCONF)
			BIT 20 	-> 	Vector Floating-Point Classification Unit (VFCLASS)
			BIT 19 	-> 	Vector Floating-Point Comparison Unit (VFCMP)
			BIT 18	-> 	Vector Floating Point Square-Root Unit (VFSQRT)
			BIT 17 	-> 	Vector Floating-Point Division Unit (VFDIV)
			BIT 16 	-> 	Vector Floating-Point Multiplication Unit (VFMUL)
			BIT 15 	-> 	Vector Floating-Point Addition Unit (VFADD)
			BIT 14 	-> 	Vector Merge Unit (VMERGE)
			BIT 13 	-> 	Vector Division Unit (VDIV)
			BIT 12 	-> 	Vector Multiplication Unit (VMUL)
			BIT 11 	-> 	Vector Comparison Unit (VCMP)
			BIT 10 	-> 	Vector Shift Unit (VSHFT)
			BIT 9 	-> 	Vector Logic Unit (VLOGIC)
			BIT 8	-> 	Vector Sign/Zero Extension Unit (VSZEXT)
			BIT 7 	-> 	Vector Add Unit (VADD)
			BIT 6 	-> 	Scalar Sign/Zero-Extension Unit (IMM)
			BIT 5 	-> 	Branch Unit (BR)
			BIT 4 	-> 	Scalar Set-On-Less-Than Unit (SLT)
			BIT 3	-> 	Scalar Shift Unit (SHFT)
			BIT 2 	-> 	Scalar Logic Unit (LOGIC)
			BIT 1 	-> 	Scalar Multiplication Unit (MUL)
			BIT 0 	-> 	Scalar Addition Unit (ADD)
			
		Register Vector
			BIT 6 	-> 	Vector v0 Register is Needed to Perform the Operation (VMASK)
			BIT 5 	-> 	Vector vs1 Register Field is Present in the Instruction Format (VS1)
			BIT 4 	-> 	Vector vs2 Register Field is Present in the Instruction Format (VS2)
			BIT 3	-> 	Vector vd Register Field is Present in the Instruction Format (VD)
			BIT 2 	-> 	Scalar rs1 Register Field is Present in the Instruction Format (RS1)
			BIT 1 	-> 	Scalar rs2 Register Field is Present in the Instruction Format (RS2)
			BIT 0 	-> 	Scalar rd Register Field is Present in the Instruction Format (RD)
			
		Operation Vector
			BIT 28 	-> 	Vector Instruction Returns the High Part of the Operation (VHL)
			BIT 27	-> 	Vector Instruction Field vs2 is Needed for Decoding (VS2)
			BIT 26	-> 	Vector Instruction Field vs1 is Needed for Decoding (VS1)
			BIT 25 	-> 	Vector Instruction Field funct6 is Needed for Decoding (F6)
			BIT 24	-> 	Vector Instruction Field vm is Needed for Decoding (VM)
			BIT 23	-> 	Vector Operand vs2's Elements are Signed (VSB)
			BIT 22	-> 	Vector Operand vs1's Elements are Signed (VSA)
			BIT 21 	-> 	Vector Memory Operation (VMEM)
			BIT 20 	-> 	Vector Fixed-Point Operation (VFXP)
			BIT 19 	-> 	Vector Floating-Point Operation (VFP)
			BIT 18	-> 	Vector Integer Operation (VINT)
			BIT 17 	-> 	Vector Operation (VEC)
			BIT 16 	-> 	Floating-Point Operation (FP)
			BIT 15 	-> 	Exception-Handling Operation (EH)
			BIT 14 	-> 	Scalar Memory Operation (MEM)
			BIT 13 	-> 	Scalar Integer Operation (INT)
			BIT 12 	-> 	opcode/funct7 is Needed for Decoding (OP/F7)
			BIT 11 	-> 	f3 is Needed for Decoding (F3)
			BIT 10 	-> 	Reserved (R)
			BIT 9 	-> 	Reserved (R)
			BIT 8	-> 	Relative-to-PC Address-Calculation Operation (PC)
			BIT 7 	-> 	Scalar rs2 is Signed (SB)
			BIT 6 	-> 	Scalar rs1 is Signed (SA)
			BIT 5 	-> 	Word's High-Part Operation (HL)
			BIT 4 	-> 	One-Word Operation (W)
			BIT 3	-> 	Atomic Memory Sync (Wait-for-Pipeline) Instruction (WP)
			BIT 2 	-> 	Conditional Branch Operation (BR)
			BIT 1 	-> 	Jump-Register Operation (JR)
			BIT 0 	-> 	Jump Operation (J)
*/
//mop
`define		unit_stride				2'b00
`define		indexed_unordered		2'b01
`define		strided					2'b10
`define		indexed_ordered			2'b11

//nf
`define		nf_1					3'b000
`define		nf_2					3'b001
`define		nf_3					3'b010
`define		nf_4					3'b011
`define		nf_5					3'b100
`define		nf_6					3'b101
`define		nf_7					3'b110
`define		nf_8					3'b111

////nf[5:3]_mew[2]_mop[1:0]
//	//LOAD
//`define		vle_w							6'b000000
//`define		vlm								6'b000000
//`define		vlse_w							6'b000010
//`define		vluxei_w						6'b000001
//`define		vloxei_w						6'b000011
//`define		vle_w_ff						6'b000000
//
//	//STORE				
//`define		vse_w							6'b000000
//`define		vsm								6'b000000
//`define		vsse_w							6'b000010
//`define		vsuxei_w						6'b000001
//`define		vsoxei_w						6'b000011
//
//	//LOAD
//`define		vlseg1e_w						6'b000000
//`define		vlseg2e_w						6'b001000
//`define		vlseg3e_w						6'b010000	
//`define		vlseg4e_w						6'b011000		
//`define		vlseg5e_w						6'b100000		
//`define		vlseg6e_w						6'b101000		
//`define		vlseg7e_w						6'b110000		
//`define		vlseg8e_w						6'b111000		
//	//STORE
//`define		vsseg1e_w						6'b000000		
//`define		vsseg2e_w						6'b001000		
//`define		vsseg3e_w						6'b010000		
//`define		vsseg4e_w						6'b011000		
//`define		vsseg5e_w						6'b100000		
//`define		vsseg6e_w						6'b101000		
//`define		vsseg7e_w						6'b110000		
//`define		vsseg8e_w						6'b111000		
//	//LOAD
//`define		vlseg1e_w_ff					6'b000000		
//`define		vlseg2e_w_ff					6'b001000		
//`define		vlseg3e_w_ff					6'b010000		
//`define		vlseg4e_w_ff					6'b011000		
//`define		vlseg5e_w_ff					6'b100000		
//`define		vlseg6e_w_ff					6'b101000		
//`define		vlseg7e_w_ff					6'b110000		
//`define		vlseg8e_w_ff					6'b111000		
//	//LOAD
//`define		vlsseg1e_w						6'b000010		
//`define		vlsseg2e_w						6'b001010		
//`define		vlsseg3e_w						6'b010010		
//`define		vlsseg4e_w						6'b011010		
//`define		vlsseg5e_w						6'b100010		
//`define		vlsseg6e_w						6'b101010		
//`define		vlsseg7e_w						6'b110010		
//`define		vlsseg8e_w						6'b111010		
//	//STORE
//`define		vssseg1e_w						6'b000010		
//`define		vssseg2e_w						6'b001010		
//`define		vssseg3e_w						6'b010010		
//`define		vssseg4e_w						6'b011010		
//`define		vssseg5e_w						6'b100010		
//`define		vssseg6e_w						6'b101010		
//`define		vssseg7e_w						6'b110010		
//`define		vssseg8e_w						6'b111010		
//	//LOAD
//`define		vluxseg1ei_w					6'b000001
//`define 	vluxseg2ei_w					6'b001001
//`define 	vluxseg3ei_w					6'b010001
//`define 	vluxseg4ei_w					6'b011001
//`define 	vluxseg5ei_w					6'b100001
//`define 	vluxseg6ei_w					6'b101001
//`define 	vluxseg7ei_w					6'b110001
//`define 	vluxseg8ei_w					6'b111001
//	//LOAD
//`define 	vloxseg1ei_w					6'b000011
//`define 	vloxseg2ei_w					6'b001011
//`define 	vloxseg3ei_w					6'b010011
//`define 	vloxseg4ei_w					6'b011011
//`define 	vloxseg5ei_w					6'b100011
//`define 	vloxseg6ei_w					6'b101011
//`define 	vloxseg7ei_w					6'b110011
//`define 	vloxseg8ei_w					6'b111011
//	//STORE
//`define 	vsuxseg1ei_w					6'b000001
//`define 	vsuxseg2ei_w					6'b001001
//`define 	vsuxseg3ei_w					6'b010001
//`define 	vsuxseg4ei_w					6'b011001
//`define 	vsuxseg5ei_w					6'b100001
//`define 	vsuxseg6ei_w					6'b101001
//`define 	vsuxseg7ei_w					6'b110001
//`define 	vsuxseg8ei_w					6'b111001
//	//STORE
//`define 	vsoxseg1ei_w					6'b000011
//`define 	vsoxseg2ei_w					6'b001011
//`define 	vsoxseg3ei_w					6'b010011
//`define 	vsoxseg4ei_w					6'b011011
//`define 	vsoxseg5ei_w					6'b100011
//`define 	vsoxseg6ei_w					6'b101011
//`define 	vsoxseg7ei_w					6'b110011
//`define 	vsoxseg8ei_w					6'b111011
//	//LOAD
//`define 	vl1re_w							6'b000000
//`define 	vl2re_w							6'b001000
//`define 	vl4re_w							6'b011000
//`define 	vl8re_w							6'b111000
//	//STORE
//`define 	vs1r							6'b000000
//`define 	vs2r							6'b001000
//`define 	vs4r							6'b011000
//`define 	vs8r							6'b111000

// funct5
`define		funct5_vle_w_ff		5'b10000

//WIDTH
`define		w8								3'b000
`define		w16								3'b101
`define		w32								3'b110
`define		w64								3'b111

//lumop_sumop	(ls=load or store, l=load)
`define		unit_stride_load_store					5'b00000
`define		unit_stride_whole_register_load_store	5'b01000
`define		unit_stride_mask_load_store				5'b01011
`define		unit_stride_fault_only_first_load		5'b10000

//data vector
	//system vector
`define 	vle8_v_system_vector				6'b000010
`define 	vle16_v_system_vector				6'b000010
`define 	vle32_v_system_vector				6'b000010
`define 	vle64_v_system_vector				6'b000010
`define 	vse8_v_system_vector				6'b000001
`define 	vse16_v_system_vector				6'b000001
`define 	vse32_v_system_vector				6'b000001
`define 	vse64_v_system_vector				6'b000001
`define 	vlm_v_system_vector					6'b000010
`define 	vsm_v_system_vector					6'b000001
`define 	vlse8_v_system_vector				6'b000010
`define 	vlse16_v_system_vector				6'b000010
`define 	vlse32_v_system_vector				6'b000010
`define 	vlse64_v_system_vector				6'b000010
`define 	vsse8_v_system_vector				6'b000001
`define 	vsse16_v_system_vector				6'b000001
`define 	vsse32_v_system_vector				6'b000001
`define 	vsse64_v_system_vector				6'b000001
`define 	vluxei8_v_system_vector				6'b000010
`define 	vluxei16_v_system_vector			6'b000010
`define 	vluxei32_v_system_vector			6'b000010
`define 	vluxei64_v_system_vector			6'b000010
`define 	vloxei8_v_system_vector				6'b000010
`define 	vloxei16_v_system_vector			6'b000010
`define 	vloxei32_v_system_vector			6'b000010
`define 	vloxei64_v_system_vector			6'b000010
`define 	vsuxei8_v_system_vector				6'b000001
`define 	vsuxei16_v_system_vector			6'b000001
`define 	vsuxei32_v_system_vector			6'b000001
`define 	vsuxei64_v_system_vector			6'b000001
`define 	vsoxei8_v_system_vector				6'b000001
`define 	vsoxei16_v_system_vector			6'b000001
`define 	vsoxei32_v_system_vector			6'b000001
`define 	vsoxei64_v_system_vector			6'b000001
`define 	vle8ff_v_system_vector				6'b000010
`define 	vle16ff_v_system_vector				6'b000010
`define 	vle32ff_v_system_vector				6'b000010
`define 	vle64ff_v_system_vector				6'b000010
`define 	vlseg1e8_v_system_vector			6'b000010
`define 	vlseg1e16_v_system_vector			6'b000010
`define 	vlseg1e32_v_system_vector			6'b000010
`define 	vlseg1e64_v_system_vector			6'b000010
`define 	vlseg2e8_v_system_vector			6'b000010
`define 	vlseg2e16_v_system_vector			6'b000010
`define 	vlseg2e32_v_system_vector			6'b000010
`define 	vlseg2e64_v_system_vector			6'b000010
`define 	vlseg3e8_v_system_vector			6'b000010
`define 	vlseg3e16_v_system_vector			6'b000010
`define 	vlseg3e32_v_system_vector			6'b000010
`define 	vlseg3e64_v_system_vector			6'b000010
`define 	vlseg4e8_v_system_vector			6'b000010
`define 	vlseg4e16_v_system_vector			6'b000010
`define 	vlseg4e32_v_system_vector			6'b000010
`define 	vlseg4e64_v_system_vector			6'b000010
`define 	vlseg5e8_v_system_vector			6'b000010
`define 	vlseg5e16_v_system_vector			6'b000010
`define 	vlseg5e32_v_system_vector			6'b000010
`define 	vlseg5e64_v_system_vector			6'b000010
`define 	vlseg6e8_v_system_vector			6'b000010
`define 	vlseg6e16_v_system_vector			6'b000010
`define 	vlseg6e32_v_system_vector			6'b000010
`define 	vlseg6e64_v_system_vector			6'b000010
`define 	vlseg7e8_v_system_vector			6'b000010
`define 	vlseg7e16_v_system_vector			6'b000010
`define 	vlseg7e32_v_system_vector			6'b000010
`define 	vlseg7e64_v_system_vector			6'b000010
`define 	vlseg8e8_v_system_vector			6'b000010
`define 	vlseg8e16_v_system_vector			6'b000010
`define 	vlseg8e32_v_system_vector			6'b000010
`define 	vlseg8e64_v_system_vector			6'b000010
`define 	vsseg1e8_v_system_vector			6'b000001
`define 	vsseg1e16_v_system_vector			6'b000001
`define 	vsseg1e32_v_system_vector			6'b000001
`define 	vsseg1e64_v_system_vector			6'b000001
`define 	vsseg2e8_v_system_vector			6'b000001
`define 	vsseg2e16_v_system_vector			6'b000001
`define 	vsseg2e32_v_system_vector			6'b000001
`define 	vsseg2e64_v_system_vector			6'b000001
`define 	vsseg3e8_v_system_vector			6'b000001
`define 	vsseg3e16_v_system_vector			6'b000001
`define 	vsseg3e32_v_system_vector			6'b000001
`define 	vsseg3e64_v_system_vector			6'b000001
`define 	vsseg4e8_v_system_vector			6'b000001
`define 	vsseg4e16_v_system_vector			6'b000001
`define 	vsseg4e32_v_system_vector			6'b000001
`define 	vsseg4e64_v_system_vector			6'b000001
`define 	vsseg5e8_v_system_vector			6'b000001
`define 	vsseg5e16_v_system_vector			6'b000001
`define 	vsseg5e32_v_system_vector			6'b000001
`define 	vsseg5e64_v_system_vector			6'b000001
`define 	vsseg6e8_v_system_vector			6'b000001
`define 	vsseg6e16_v_system_vector			6'b000001
`define 	vsseg6e32_v_system_vector			6'b000001
`define 	vsseg6e64_v_system_vector			6'b000001
`define 	vsseg7e8_v_system_vector			6'b000001
`define 	vsseg7e16_v_system_vector			6'b000001
`define 	vsseg7e32_v_system_vector			6'b000001
`define 	vsseg7e64_v_system_vector			6'b000001
`define 	vsseg8e8_v_system_vector			6'b000001
`define 	vsseg8e16_v_system_vector			6'b000001
`define 	vsseg8e32_v_system_vector			6'b000001
`define 	vsseg8e64_v_system_vector			6'b000001
`define 	vlseg1e8ff_v_system_vector			6'b000010
`define 	vlseg1e16ff_v_system_vector			6'b000010
`define 	vlseg1e32ff_v_system_vector			6'b000010
`define 	vlseg1e64ff_v_system_vector			6'b000010
`define 	vlseg2e8ff_v_system_vector			6'b000010
`define 	vlseg2e16ff_v_system_vector			6'b000010
`define 	vlseg2e32ff_v_system_vector			6'b000010
`define 	vlseg2e64ff_v_system_vector			6'b000010
`define 	vlseg3e8ff_v_system_vector			6'b000010
`define 	vlseg3e16ff_v_system_vector			6'b000010
`define 	vlseg3e32ff_v_system_vector			6'b000010
`define 	vlseg3e64ff_v_system_vector			6'b000010
`define 	vlseg4e8ff_v_system_vector			6'b000010
`define 	vlseg4e16ff_v_system_vector			6'b000010
`define 	vlseg4e32ff_v_system_vector			6'b000010
`define 	vlseg4e64ff_v_system_vector			6'b000010
`define 	vlseg5e8ff_v_system_vector			6'b000010
`define 	vlseg5e16ff_v_system_vector			6'b000010
`define 	vlseg5e32ff_v_system_vector			6'b000010
`define 	vlseg5e64ff_v_system_vector			6'b000010
`define 	vlseg6e8ff_v_system_vector			6'b000010
`define 	vlseg6e16ff_v_system_vector			6'b000010
`define 	vlseg6e32ff_v_system_vector			6'b000010
`define 	vlseg6e64ff_v_system_vector			6'b000010
`define 	vlseg7e8ff_v_system_vector			6'b000010
`define 	vlseg7e16ff_v_system_vector			6'b000010
`define 	vlseg7e32ff_v_system_vector			6'b000010
`define 	vlseg7e64ff_v_system_vector			6'b000010
`define 	vlseg8e8ff_v_system_vector			6'b000010
`define 	vlseg8e16ff_v_system_vector			6'b000010
`define 	vlseg8e32ff_v_system_vector			6'b000010
`define 	vlseg8e64ff_v_system_vector			6'b000010
`define 	vlsseg1e8_v_system_vector			6'b000010
`define 	vlsseg1e16_v_system_vector			6'b000010
`define 	vlsseg1e32_v_system_vector			6'b000010
`define 	vlsseg1e64_v_system_vector			6'b000010
`define 	vlsseg2e8_v_system_vector			6'b000010
`define 	vlsseg2e16_v_system_vector			6'b000010
`define 	vlsseg2e32_v_system_vector			6'b000010
`define 	vlsseg2e64_v_system_vector			6'b000010
`define 	vlsseg3e8_v_system_vector			6'b000010
`define 	vlsseg3e16_v_system_vector			6'b000010
`define 	vlsseg3e32_v_system_vector			6'b000010
`define 	vlsseg3e64_v_system_vector			6'b000010
`define 	vlsseg4e8_v_system_vector			6'b000010
`define 	vlsseg4e16_v_system_vector			6'b000010
`define 	vlsseg4e32_v_system_vector			6'b000010
`define 	vlsseg4e64_v_system_vector			6'b000010
`define 	vlsseg5e8_v_system_vector			6'b000010
`define 	vlsseg5e16_v_system_vector			6'b000010
`define 	vlsseg5e32_v_system_vector			6'b000010
`define 	vlsseg5e64_v_system_vector			6'b000010
`define 	vlsseg6e8_v_system_vector			6'b000010
`define 	vlsseg6e16_v_system_vector			6'b000010
`define 	vlsseg6e32_v_system_vector			6'b000010
`define 	vlsseg6e64_v_system_vector			6'b000010
`define 	vlsseg7e8_v_system_vector			6'b000010
`define 	vlsseg7e16_v_system_vector			6'b000010
`define 	vlsseg7e32_v_system_vector			6'b000010
`define 	vlsseg7e64_v_system_vector			6'b000010
`define 	vlsseg8e8_v_system_vector			6'b000010
`define 	vlsseg8e16_v_system_vector			6'b000010
`define 	vlsseg8e32_v_system_vector			6'b000010
`define 	vlsseg8e64_v_system_vector			6'b000010
`define 	vssseg1e8_v_system_vector			6'b000001
`define 	vssseg1e16_v_system_vector			6'b000001
`define 	vssseg1e32_v_system_vector			6'b000001
`define 	vssseg1e64_v_system_vector			6'b000001
`define 	vssseg2e8_v_system_vector			6'b000001
`define 	vssseg2e16_v_system_vector			6'b000001
`define 	vssseg2e32_v_system_vector			6'b000001
`define 	vssseg2e64_v_system_vector			6'b000001
`define 	vssseg3e8_v_system_vector			6'b000001
`define 	vssseg3e16_v_system_vector			6'b000001
`define 	vssseg3e32_v_system_vector			6'b000001
`define 	vssseg3e64_v_system_vector			6'b000001
`define 	vssseg4e8_v_system_vector			6'b000001
`define 	vssseg4e16_v_system_vector			6'b000001
`define 	vssseg4e32_v_system_vector			6'b000001
`define 	vssseg4e64_v_system_vector			6'b000001
`define 	vssseg5e8_v_system_vector			6'b000001
`define 	vssseg5e16_v_system_vector			6'b000001
`define 	vssseg5e32_v_system_vector			6'b000001
`define 	vssseg5e64_v_system_vector			6'b000001
`define 	vssseg6e8_v_system_vector			6'b000001
`define 	vssseg6e16_v_system_vector			6'b000001
`define 	vssseg6e32_v_system_vector			6'b000001
`define 	vssseg6e64_v_system_vector			6'b000001
`define 	vssseg7e8_v_system_vector			6'b000001
`define 	vssseg7e16_v_system_vector			6'b000001
`define 	vssseg7e32_v_system_vector			6'b000001
`define 	vssseg7e64_v_system_vector			6'b000001
`define 	vssseg8e8_v_system_vector			6'b000001
`define 	vssseg8e16_v_system_vector			6'b000001
`define 	vssseg8e32_v_system_vector			6'b000001
`define 	vssseg8e64_v_system_vector			6'b000001
`define 	vluxseg1ei8_v_system_vector			6'b000010
`define 	vluxseg1ei16_v_system_vector		6'b000010
`define 	vluxseg1ei32_v_system_vector		6'b000010
`define 	vluxseg1ei64_v_system_vector		6'b000010
`define 	vluxseg2ei8_v_system_vector			6'b000010
`define 	vluxseg2ei16_v_system_vector		6'b000010
`define 	vluxseg2ei32_v_system_vector		6'b000010
`define 	vluxseg2ei64_v_system_vector		6'b000010
`define 	vluxseg3ei8_v_system_vector			6'b000010
`define 	vluxseg3ei16_v_system_vector		6'b000010
`define 	vluxseg3ei32_v_system_vector		6'b000010
`define 	vluxseg3ei64_v_system_vector		6'b000010
`define 	vluxseg4ei8_v_system_vector			6'b000010
`define 	vluxseg4ei16_v_system_vector		6'b000010
`define 	vluxseg4ei32_v_system_vector		6'b000010
`define 	vluxseg4ei64_v_system_vector		6'b000010
`define 	vluxseg5ei8_v_system_vector			6'b000010
`define 	vluxseg5ei16_v_system_vector		6'b000010
`define 	vluxseg5ei32_v_system_vector		6'b000010
`define 	vluxseg5ei64_v_system_vector		6'b000010
`define 	vluxseg6ei8_v_system_vector			6'b000010
`define 	vluxseg6ei16_v_system_vector		6'b000010
`define 	vluxseg6ei32_v_system_vector		6'b000010
`define 	vluxseg6ei64_v_system_vector		6'b000010
`define 	vluxseg7ei8_v_system_vector			6'b000010
`define 	vluxseg7ei16_v_system_vector		6'b000010
`define 	vluxseg7ei32_v_system_vector		6'b000010
`define 	vluxseg7ei64_v_system_vector		6'b000010
`define 	vluxseg8ei8_v_system_vector			6'b000010
`define 	vluxseg8ei16_v_system_vector		6'b000010
`define 	vluxseg8ei32_v_system_vector		6'b000010
`define 	vluxseg8ei64_v_system_vector		6'b000010
`define 	vloxseg1ei8_v_system_vector			6'b000010
`define 	vloxseg1ei16_v_system_vector		6'b000010
`define 	vloxseg1ei32_v_system_vector		6'b000010
`define 	vloxseg1ei64_v_system_vector		6'b000010
`define 	vloxseg2ei8_v_system_vector			6'b000010
`define 	vloxseg2ei16_v_system_vector		6'b000010
`define 	vloxseg2ei32_v_system_vector		6'b000010
`define 	vloxseg2ei64_v_system_vector		6'b000010
`define 	vloxseg3ei8_v_system_vector			6'b000010
`define 	vloxseg3ei16_v_system_vector		6'b000010
`define 	vloxseg3ei32_v_system_vector		6'b000010
`define 	vloxseg3ei64_v_system_vector		6'b000010
`define 	vloxseg4ei8_v_system_vector			6'b000010
`define 	vloxseg4ei16_v_system_vector		6'b000010
`define 	vloxseg4ei32_v_system_vector		6'b000010
`define 	vloxseg4ei64_v_system_vector		6'b000010
`define 	vloxseg5ei8_v_system_vector			6'b000010
`define 	vloxseg5ei16_v_system_vector		6'b000010
`define 	vloxseg5ei32_v_system_vector		6'b000010
`define 	vloxseg5ei64_v_system_vector		6'b000010
`define 	vloxseg6ei8_v_system_vector			6'b000010
`define 	vloxseg6ei16_v_system_vector		6'b000010
`define 	vloxseg6ei32_v_system_vector		6'b000010
`define 	vloxseg6ei64_v_system_vector		6'b000010
`define 	vloxseg7ei8_v_system_vector			6'b000010
`define 	vloxseg7ei16_v_system_vector		6'b000010
`define 	vloxseg7ei32_v_system_vector		6'b000010
`define 	vloxseg7ei64_v_system_vector		6'b000010
`define 	vloxseg8ei8_v_system_vector			6'b000010
`define 	vloxseg8ei16_v_system_vector		6'b000010
`define 	vloxseg8ei32_v_system_vector		6'b000010
`define 	vloxseg8ei64_v_system_vector		6'b000010
`define 	vsuxseg1ei8_v_system_vector			6'b000001
`define 	vsuxseg1ei16_v_system_vector		6'b000001
`define 	vsuxseg1ei32_v_system_vector		6'b000001
`define 	vsuxseg1ei64_v_system_vector		6'b000001
`define 	vsuxseg2ei8_v_system_vector			6'b000001
`define 	vsuxseg2ei16_v_system_vector		6'b000001
`define 	vsuxseg2ei32_v_system_vector		6'b000001
`define 	vsuxseg2ei64_v_system_vector		6'b000001
`define 	vsuxseg3ei8_v_system_vector			6'b000001
`define 	vsuxseg3ei16_v_system_vector		6'b000001
`define 	vsuxseg3ei32_v_system_vector		6'b000001
`define 	vsuxseg3ei64_v_system_vector		6'b000001
`define 	vsuxseg4ei8_v_system_vector			6'b000001
`define 	vsuxseg4ei16_v_system_vector		6'b000001
`define 	vsuxseg4ei32_v_system_vector		6'b000001
`define 	vsuxseg4ei64_v_system_vector		6'b000001
`define 	vsuxseg5ei8_v_system_vector			6'b000001
`define 	vsuxseg5ei16_v_system_vector		6'b000001
`define 	vsuxseg5ei32_v_system_vector		6'b000001
`define 	vsuxseg5ei64_v_system_vector		6'b000001
`define 	vsuxseg6ei8_v_system_vector			6'b000001
`define 	vsuxseg6ei16_v_system_vector		6'b000001
`define 	vsuxseg6ei32_v_system_vector		6'b000001
`define 	vsuxseg6ei64_v_system_vector		6'b000001
`define 	vsuxseg7ei8_v_system_vector			6'b000001
`define 	vsuxseg7ei16_v_system_vector		6'b000001
`define 	vsuxseg7ei32_v_system_vector		6'b000001
`define 	vsuxseg7ei64_v_system_vector		6'b000001
`define 	vsuxseg8ei8_v_system_vector			6'b000001
`define 	vsuxseg8ei16_v_system_vector		6'b000001
`define 	vsuxseg8ei32_v_system_vector		6'b000001
`define 	vsuxseg8ei64_v_system_vector		6'b000001
`define 	vsoxseg1ei8_v_system_vector			6'b000001
`define 	vsoxseg1ei16_v_system_vector		6'b000001
`define 	vsoxseg1ei32_v_system_vector		6'b000001
`define 	vsoxseg1ei64_v_system_vector		6'b000001
`define 	vsoxseg2ei8_v_system_vector			6'b000001
`define 	vsoxseg2ei16_v_system_vector		6'b000001
`define 	vsoxseg2ei32_v_system_vector		6'b000001
`define 	vsoxseg2ei64_v_system_vector		6'b000001
`define 	vsoxseg3ei8_v_system_vector			6'b000001
`define 	vsoxseg3ei16_v_system_vector		6'b000001
`define 	vsoxseg3ei32_v_system_vector		6'b000001
`define 	vsoxseg3ei64_v_system_vector		6'b000001
`define 	vsoxseg4ei8_v_system_vector			6'b000001
`define 	vsoxseg4ei16_v_system_vector		6'b000001
`define 	vsoxseg4ei32_v_system_vector		6'b000001
`define 	vsoxseg4ei64_v_system_vector		6'b000001
`define 	vsoxseg5ei8_v_system_vector			6'b000001
`define 	vsoxseg5ei16_v_system_vector		6'b000001
`define 	vsoxseg5ei32_v_system_vector		6'b000001
`define 	vsoxseg5ei64_v_system_vector		6'b000001
`define 	vsoxseg6ei8_v_system_vector			6'b000001
`define 	vsoxseg6ei16_v_system_vector		6'b000001
`define 	vsoxseg6ei32_v_system_vector		6'b000001
`define 	vsoxseg6ei64_v_system_vector		6'b000001
`define 	vsoxseg7ei8_v_system_vector			6'b000001
`define 	vsoxseg7ei16_v_system_vector		6'b000001
`define 	vsoxseg7ei32_v_system_vector		6'b000001
`define 	vsoxseg7ei64_v_system_vector		6'b000001
`define 	vsoxseg8ei8_v_system_vector			6'b000001
`define 	vsoxseg8ei16_v_system_vector		6'b000001
`define 	vsoxseg8ei32_v_system_vector		6'b000001
`define 	vsoxseg8ei64_v_system_vector		6'b000001
`define 	vl1re8_v_system_vector				6'b000010
`define 	vl1re16_v_system_vector				6'b000010
`define 	vl1re32_v_system_vector				6'b000010
`define 	vl1re64_v_system_vector				6'b000010
`define 	vl2re8_v_system_vector				6'b000010
`define 	vl2re16_v_system_vector				6'b000010
`define 	vl2re32_v_system_vector				6'b000010
`define 	vl2re64_v_system_vector				6'b000010
`define 	vl4re8_v_system_vector				6'b000010
`define 	vl4re16_v_system_vector				6'b000010
`define 	vl4re32_v_system_vector				6'b000010
`define 	vl4re64_v_system_vector				6'b000010
`define 	vl8re8_v_system_vector				6'b000010
`define 	vl8re16_v_system_vector				6'b000010
`define 	vl8re32_v_system_vector				6'b000010
`define 	vl8re64_v_system_vector				6'b000010
`define 	vs1r_v_system_vector				6'b000001
`define 	vs2r_v_system_vector				6'b000001
`define 	vs4r_v_system_vector				6'b000001
`define 	vs8r_v_system_vector				6'b000001

	//resource vector
`define 	vle8_v_resource_vector				22'b0000000000000000000000
`define 	vle16_v_resource_vector				22'b0000000000000000000000
`define 	vle32_v_resource_vector				22'b0000000000000000000000
`define 	vle64_v_resource_vector				22'b0000000000000000000000
`define 	vse8_v_resource_vector				22'b0000000000000000000000
`define 	vse16_v_resource_vector				22'b0000000000000000000000
`define 	vse32_v_resource_vector				22'b0000000000000000000000
`define 	vse64_v_resource_vector				22'b0000000000000000000000
`define 	vlm_v_resource_vector				22'b0000000000000000000000
`define 	vsm_v_resource_vector				22'b0000000000000000000000
`define 	vlse8_v_resource_vector				22'b0000000000000000000000
`define 	vlse16_v_resource_vector			22'b0000000000000000000000
`define 	vlse32_v_resource_vector			22'b0000000000000000000000
`define 	vlse64_v_resource_vector			22'b0000000000000000000000
`define 	vsse8_v_resource_vector				22'b0000000000000000000000
`define 	vsse16_v_resource_vector			22'b0000000000000000000000
`define 	vsse32_v_resource_vector			22'b0000000000000000000000
`define 	vsse64_v_resource_vector			22'b0000000000000000000000
`define 	vluxei8_v_resource_vector			22'b0000000000000000000000
`define 	vluxei16_v_resource_vector			22'b0000000000000000000000
`define 	vluxei32_v_resource_vector			22'b0000000000000000000000
`define 	vluxei64_v_resource_vector			22'b0000000000000000000000
`define 	vloxei8_v_resource_vector			22'b0000000000000000000000
`define 	vloxei16_v_resource_vector			22'b0000000000000000000000
`define 	vloxei32_v_resource_vector			22'b0000000000000000000000
`define 	vloxei64_v_resource_vector			22'b0000000000000000000000
`define 	vsuxei8_v_resource_vector			22'b0000000000000000000000
`define 	vsuxei16_v_resource_vector			22'b0000000000000000000000
`define 	vsuxei32_v_resource_vector			22'b0000000000000000000000
`define 	vsuxei64_v_resource_vector			22'b0000000000000000000000
`define 	vsoxei8_v_resource_vector			22'b0000000000000000000000
`define 	vsoxei16_v_resource_vector			22'b0000000000000000000000
`define 	vsoxei32_v_resource_vector			22'b0000000000000000000000
`define 	vsoxei64_v_resource_vector			22'b0000000000000000000000
`define 	vle8ff_v_resource_vector			22'b0000000000000000000000
`define 	vle16ff_v_resource_vector			22'b0000000000000000000000
`define 	vle32ff_v_resource_vector			22'b0000000000000000000000
`define 	vle64ff_v_resource_vector			22'b0000000000000000000000
`define 	vlseg1e8_v_resource_vector			22'b0000000000000000000000
`define 	vlseg1e16_v_resource_vector			22'b0000000000000000000000
`define 	vlseg1e32_v_resource_vector			22'b0000000000000000000000
`define 	vlseg1e64_v_resource_vector			22'b0000000000000000000000
`define 	vlseg2e8_v_resource_vector			22'b0000000000000000000000
`define 	vlseg2e16_v_resource_vector			22'b0000000000000000000000
`define 	vlseg2e32_v_resource_vector			22'b0000000000000000000000
`define 	vlseg2e64_v_resource_vector			22'b0000000000000000000000
`define 	vlseg3e8_v_resource_vector			22'b0000000000000000000000
`define 	vlseg3e16_v_resource_vector			22'b0000000000000000000000
`define 	vlseg3e32_v_resource_vector			22'b0000000000000000000000
`define 	vlseg3e64_v_resource_vector			22'b0000000000000000000000
`define 	vlseg4e8_v_resource_vector			22'b0000000000000000000000
`define 	vlseg4e16_v_resource_vector			22'b0000000000000000000000
`define 	vlseg4e32_v_resource_vector			22'b0000000000000000000000
`define 	vlseg4e64_v_resource_vector			22'b0000000000000000000000
`define 	vlseg5e8_v_resource_vector			22'b0000000000000000000000
`define 	vlseg5e16_v_resource_vector			22'b0000000000000000000000
`define 	vlseg5e32_v_resource_vector			22'b0000000000000000000000
`define 	vlseg5e64_v_resource_vector			22'b0000000000000000000000
`define 	vlseg6e8_v_resource_vector			22'b0000000000000000000000
`define 	vlseg6e16_v_resource_vector			22'b0000000000000000000000
`define 	vlseg6e32_v_resource_vector			22'b0000000000000000000000
`define 	vlseg6e64_v_resource_vector			22'b0000000000000000000000
`define 	vlseg7e8_v_resource_vector			22'b0000000000000000000000
`define 	vlseg7e16_v_resource_vector			22'b0000000000000000000000
`define 	vlseg7e32_v_resource_vector			22'b0000000000000000000000
`define 	vlseg7e64_v_resource_vector			22'b0000000000000000000000
`define 	vlseg8e8_v_resource_vector			22'b0000000000000000000000
`define 	vlseg8e16_v_resource_vector			22'b0000000000000000000000
`define 	vlseg8e32_v_resource_vector			22'b0000000000000000000000
`define 	vlseg8e64_v_resource_vector			22'b0000000000000000000000
`define 	vsseg1e8_v_resource_vector			22'b0000000000000000000000
`define 	vsseg1e16_v_resource_vector			22'b0000000000000000000000
`define 	vsseg1e32_v_resource_vector			22'b0000000000000000000000
`define 	vsseg1e64_v_resource_vector			22'b0000000000000000000000
`define 	vsseg2e8_v_resource_vector			22'b0000000000000000000000
`define 	vsseg2e16_v_resource_vector			22'b0000000000000000000000
`define 	vsseg2e32_v_resource_vector			22'b0000000000000000000000
`define 	vsseg2e64_v_resource_vector			22'b0000000000000000000000
`define 	vsseg3e8_v_resource_vector			22'b0000000000000000000000
`define 	vsseg3e16_v_resource_vector			22'b0000000000000000000000
`define 	vsseg3e32_v_resource_vector			22'b0000000000000000000000
`define 	vsseg3e64_v_resource_vector			22'b0000000000000000000000
`define 	vsseg4e8_v_resource_vector			22'b0000000000000000000000
`define 	vsseg4e16_v_resource_vector			22'b0000000000000000000000
`define 	vsseg4e32_v_resource_vector			22'b0000000000000000000000
`define 	vsseg4e64_v_resource_vector			22'b0000000000000000000000
`define 	vsseg5e8_v_resource_vector			22'b0000000000000000000000
`define 	vsseg5e16_v_resource_vector			22'b0000000000000000000000
`define 	vsseg5e32_v_resource_vector			22'b0000000000000000000000
`define 	vsseg5e64_v_resource_vector			22'b0000000000000000000000
`define 	vsseg6e8_v_resource_vector			22'b0000000000000000000000
`define 	vsseg6e16_v_resource_vector			22'b0000000000000000000000
`define 	vsseg6e32_v_resource_vector			22'b0000000000000000000000
`define 	vsseg6e64_v_resource_vector			22'b0000000000000000000000
`define 	vsseg7e8_v_resource_vector			22'b0000000000000000000000
`define 	vsseg7e16_v_resource_vector			22'b0000000000000000000000
`define 	vsseg7e32_v_resource_vector			22'b0000000000000000000000
`define 	vsseg7e64_v_resource_vector			22'b0000000000000000000000
`define 	vsseg8e8_v_resource_vector			22'b0000000000000000000000
`define 	vsseg8e16_v_resource_vector			22'b0000000000000000000000
`define 	vsseg8e32_v_resource_vector			22'b0000000000000000000000
`define 	vsseg8e64_v_resource_vector			22'b0000000000000000000000
`define 	vlseg1e8ff_v_resource_vector		22'b0000000000000000000000
`define 	vlseg1e16ff_v_resource_vector		22'b0000000000000000000000
`define 	vlseg1e32ff_v_resource_vector		22'b0000000000000000000000
`define 	vlseg1e64ff_v_resource_vector		22'b0000000000000000000000
`define 	vlseg2e8ff_v_resource_vector		22'b0000000000000000000000
`define 	vlseg2e16ff_v_resource_vector		22'b0000000000000000000000
`define 	vlseg2e32ff_v_resource_vector		22'b0000000000000000000000
`define 	vlseg2e64ff_v_resource_vector		22'b0000000000000000000000
`define 	vlseg3e8ff_v_resource_vector		22'b0000000000000000000000
`define 	vlseg3e16ff_v_resource_vector		22'b0000000000000000000000
`define 	vlseg3e32ff_v_resource_vector		22'b0000000000000000000000
`define 	vlseg3e64ff_v_resource_vector		22'b0000000000000000000000
`define 	vlseg4e8ff_v_resource_vector		22'b0000000000000000000000
`define 	vlseg4e16ff_v_resource_vector		22'b0000000000000000000000
`define 	vlseg4e32ff_v_resource_vector		22'b0000000000000000000000
`define 	vlseg4e64ff_v_resource_vector		22'b0000000000000000000000
`define 	vlseg5e8ff_v_resource_vector		22'b0000000000000000000000
`define 	vlseg5e16ff_v_resource_vector		22'b0000000000000000000000
`define 	vlseg5e32ff_v_resource_vector		22'b0000000000000000000000
`define 	vlseg5e64ff_v_resource_vector		22'b0000000000000000000000
`define 	vlseg6e8ff_v_resource_vector		22'b0000000000000000000000
`define 	vlseg6e16ff_v_resource_vector		22'b0000000000000000000000
`define 	vlseg6e32ff_v_resource_vector		22'b0000000000000000000000
`define 	vlseg6e64ff_v_resource_vector		22'b0000000000000000000000
`define 	vlseg7e8ff_v_resource_vector		22'b0000000000000000000000
`define 	vlseg7e16ff_v_resource_vector		22'b0000000000000000000000
`define 	vlseg7e32ff_v_resource_vector		22'b0000000000000000000000
`define 	vlseg7e64ff_v_resource_vector		22'b0000000000000000000000
`define 	vlseg8e8ff_v_resource_vector		22'b0000000000000000000000
`define 	vlseg8e16ff_v_resource_vector		22'b0000000000000000000000
`define 	vlseg8e32ff_v_resource_vector		22'b0000000000000000000000
`define 	vlseg8e64ff_v_resource_vector		22'b0000000000000000000000
`define 	vlsseg1e8_v_resource_vector			22'b0000000000000000000000
`define 	vlsseg1e16_v_resource_vector		22'b0000000000000000000000
`define 	vlsseg1e32_v_resource_vector		22'b0000000000000000000000
`define 	vlsseg1e64_v_resource_vector		22'b0000000000000000000000
`define 	vlsseg2e8_v_resource_vector			22'b0000000000000000000000
`define 	vlsseg2e16_v_resource_vector		22'b0000000000000000000000
`define 	vlsseg2e32_v_resource_vector		22'b0000000000000000000000
`define 	vlsseg2e64_v_resource_vector		22'b0000000000000000000000
`define 	vlsseg3e8_v_resource_vector			22'b0000000000000000000000
`define 	vlsseg3e16_v_resource_vector		22'b0000000000000000000000
`define 	vlsseg3e32_v_resource_vector		22'b0000000000000000000000
`define 	vlsseg3e64_v_resource_vector		22'b0000000000000000000000
`define 	vlsseg4e8_v_resource_vector			22'b0000000000000000000000
`define 	vlsseg4e16_v_resource_vector		22'b0000000000000000000000
`define 	vlsseg4e32_v_resource_vector		22'b0000000000000000000000
`define 	vlsseg4e64_v_resource_vector		22'b0000000000000000000000
`define 	vlsseg5e8_v_resource_vector			22'b0000000000000000000000
`define 	vlsseg5e16_v_resource_vector		22'b0000000000000000000000
`define 	vlsseg5e32_v_resource_vector		22'b0000000000000000000000
`define 	vlsseg5e64_v_resource_vector		22'b0000000000000000000000
`define 	vlsseg6e8_v_resource_vector			22'b0000000000000000000000
`define 	vlsseg6e16_v_resource_vector		22'b0000000000000000000000
`define 	vlsseg6e32_v_resource_vector		22'b0000000000000000000000
`define 	vlsseg6e64_v_resource_vector		22'b0000000000000000000000
`define 	vlsseg7e8_v_resource_vector			22'b0000000000000000000000
`define 	vlsseg7e16_v_resource_vector		22'b0000000000000000000000
`define 	vlsseg7e32_v_resource_vector		22'b0000000000000000000000
`define 	vlsseg7e64_v_resource_vector		22'b0000000000000000000000
`define 	vlsseg8e8_v_resource_vector			22'b0000000000000000000000
`define 	vlsseg8e16_v_resource_vector		22'b0000000000000000000000
`define 	vlsseg8e32_v_resource_vector		22'b0000000000000000000000
`define 	vlsseg8e64_v_resource_vector		22'b0000000000000000000000
`define 	vssseg1e8_v_resource_vector			22'b0000000000000000000000
`define 	vssseg1e16_v_resource_vector		22'b0000000000000000000000
`define 	vssseg1e32_v_resource_vector		22'b0000000000000000000000
`define 	vssseg1e64_v_resource_vector		22'b0000000000000000000000
`define 	vssseg2e8_v_resource_vector			22'b0000000000000000000000
`define 	vssseg2e16_v_resource_vector		22'b0000000000000000000000
`define 	vssseg2e32_v_resource_vector		22'b0000000000000000000000
`define 	vssseg2e64_v_resource_vector		22'b0000000000000000000000
`define 	vssseg3e8_v_resource_vector			22'b0000000000000000000000
`define 	vssseg3e16_v_resource_vector		22'b0000000000000000000000
`define 	vssseg3e32_v_resource_vector		22'b0000000000000000000000
`define 	vssseg3e64_v_resource_vector		22'b0000000000000000000000
`define 	vssseg4e8_v_resource_vector			22'b0000000000000000000000
`define 	vssseg4e16_v_resource_vector		22'b0000000000000000000000
`define 	vssseg4e32_v_resource_vector		22'b0000000000000000000000
`define 	vssseg4e64_v_resource_vector		22'b0000000000000000000000
`define 	vssseg5e8_v_resource_vector			22'b0000000000000000000000
`define 	vssseg5e16_v_resource_vector		22'b0000000000000000000000
`define 	vssseg5e32_v_resource_vector		22'b0000000000000000000000
`define 	vssseg5e64_v_resource_vector		22'b0000000000000000000000
`define 	vssseg6e8_v_resource_vector			22'b0000000000000000000000
`define 	vssseg6e16_v_resource_vector		22'b0000000000000000000000
`define 	vssseg6e32_v_resource_vector		22'b0000000000000000000000
`define 	vssseg6e64_v_resource_vector		22'b0000000000000000000000
`define 	vssseg7e8_v_resource_vector			22'b0000000000000000000000
`define 	vssseg7e16_v_resource_vector		22'b0000000000000000000000
`define 	vssseg7e32_v_resource_vector		22'b0000000000000000000000
`define 	vssseg7e64_v_resource_vector		22'b0000000000000000000000
`define 	vssseg8e8_v_resource_vector			22'b0000000000000000000000
`define 	vssseg8e16_v_resource_vector		22'b0000000000000000000000
`define 	vssseg8e32_v_resource_vector		22'b0000000000000000000000
`define 	vssseg8e64_v_resource_vector		22'b0000000000000000000000
`define 	vluxseg1ei8_v_resource_vector		22'b0000000000000000000000
`define 	vluxseg1ei16_v_resource_vector		22'b0000000000000000000000
`define 	vluxseg1ei32_v_resource_vector		22'b0000000000000000000000
`define 	vluxseg1ei64_v_resource_vector		22'b0000000000000000000000
`define 	vluxseg2ei8_v_resource_vector		22'b0000000000000000000000
`define 	vluxseg2ei16_v_resource_vector		22'b0000000000000000000000
`define 	vluxseg2ei32_v_resource_vector		22'b0000000000000000000000
`define 	vluxseg2ei64_v_resource_vector		22'b0000000000000000000000
`define 	vluxseg3ei8_v_resource_vector		22'b0000000000000000000000
`define 	vluxseg3ei16_v_resource_vector		22'b0000000000000000000000
`define 	vluxseg3ei32_v_resource_vector		22'b0000000000000000000000
`define 	vluxseg3ei64_v_resource_vector		22'b0000000000000000000000
`define 	vluxseg4ei8_v_resource_vector		22'b0000000000000000000000
`define 	vluxseg4ei16_v_resource_vector		22'b0000000000000000000000
`define 	vluxseg4ei32_v_resource_vector		22'b0000000000000000000000
`define 	vluxseg4ei64_v_resource_vector		22'b0000000000000000000000
`define 	vluxseg5ei8_v_resource_vector		22'b0000000000000000000000
`define 	vluxseg5ei16_v_resource_vector		22'b0000000000000000000000
`define 	vluxseg5ei32_v_resource_vector		22'b0000000000000000000000
`define 	vluxseg5ei64_v_resource_vector		22'b0000000000000000000000
`define 	vluxseg6ei8_v_resource_vector		22'b0000000000000000000000
`define 	vluxseg6ei16_v_resource_vector		22'b0000000000000000000000
`define 	vluxseg6ei32_v_resource_vector		22'b0000000000000000000000
`define 	vluxseg6ei64_v_resource_vector		22'b0000000000000000000000
`define 	vluxseg7ei8_v_resource_vector		22'b0000000000000000000000
`define 	vluxseg7ei16_v_resource_vector		22'b0000000000000000000000
`define 	vluxseg7ei32_v_resource_vector		22'b0000000000000000000000
`define 	vluxseg7ei64_v_resource_vector		22'b0000000000000000000000
`define 	vluxseg8ei8_v_resource_vector		22'b0000000000000000000000
`define 	vluxseg8ei16_v_resource_vector		22'b0000000000000000000000
`define 	vluxseg8ei32_v_resource_vector		22'b0000000000000000000000
`define 	vluxseg8ei64_v_resource_vector		22'b0000000000000000000000
`define 	vloxseg1ei8_v_resource_vector		22'b0000000000000000000000
`define 	vloxseg1ei16_v_resource_vector		22'b0000000000000000000000
`define 	vloxseg1ei32_v_resource_vector		22'b0000000000000000000000
`define 	vloxseg1ei64_v_resource_vector		22'b0000000000000000000000
`define 	vloxseg2ei8_v_resource_vector		22'b0000000000000000000000
`define 	vloxseg2ei16_v_resource_vector		22'b0000000000000000000000
`define 	vloxseg2ei32_v_resource_vector		22'b0000000000000000000000
`define 	vloxseg2ei64_v_resource_vector		22'b0000000000000000000000
`define 	vloxseg3ei8_v_resource_vector		22'b0000000000000000000000
`define 	vloxseg3ei16_v_resource_vector		22'b0000000000000000000000
`define 	vloxseg3ei32_v_resource_vector		22'b0000000000000000000000
`define 	vloxseg3ei64_v_resource_vector		22'b0000000000000000000000
`define 	vloxseg4ei8_v_resource_vector		22'b0000000000000000000000
`define 	vloxseg4ei16_v_resource_vector		22'b0000000000000000000000
`define 	vloxseg4ei32_v_resource_vector		22'b0000000000000000000000
`define 	vloxseg4ei64_v_resource_vector		22'b0000000000000000000000
`define 	vloxseg5ei8_v_resource_vector		22'b0000000000000000000000
`define 	vloxseg5ei16_v_resource_vector		22'b0000000000000000000000
`define 	vloxseg5ei32_v_resource_vector		22'b0000000000000000000000
`define 	vloxseg5ei64_v_resource_vector		22'b0000000000000000000000
`define 	vloxseg6ei8_v_resource_vector		22'b0000000000000000000000
`define 	vloxseg6ei16_v_resource_vector		22'b0000000000000000000000
`define 	vloxseg6ei32_v_resource_vector		22'b0000000000000000000000
`define 	vloxseg6ei64_v_resource_vector		22'b0000000000000000000000
`define 	vloxseg7ei8_v_resource_vector		22'b0000000000000000000000
`define 	vloxseg7ei16_v_resource_vector		22'b0000000000000000000000
`define 	vloxseg7ei32_v_resource_vector		22'b0000000000000000000000
`define 	vloxseg7ei64_v_resource_vector		22'b0000000000000000000000
`define 	vloxseg8ei8_v_resource_vector		22'b0000000000000000000000
`define 	vloxseg8ei16_v_resource_vector		22'b0000000000000000000000
`define 	vloxseg8ei32_v_resource_vector		22'b0000000000000000000000
`define 	vloxseg8ei64_v_resource_vector		22'b0000000000000000000000
`define 	vsuxseg1ei8_v_resource_vector		22'b0000000000000000000000
`define 	vsuxseg1ei16_v_resource_vector		22'b0000000000000000000000
`define 	vsuxseg1ei32_v_resource_vector		22'b0000000000000000000000
`define 	vsuxseg1ei64_v_resource_vector		22'b0000000000000000000000
`define 	vsuxseg2ei8_v_resource_vector		22'b0000000000000000000000
`define 	vsuxseg2ei16_v_resource_vector		22'b0000000000000000000000
`define 	vsuxseg2ei32_v_resource_vector		22'b0000000000000000000000
`define 	vsuxseg2ei64_v_resource_vector		22'b0000000000000000000000
`define 	vsuxseg3ei8_v_resource_vector		22'b0000000000000000000000
`define 	vsuxseg3ei16_v_resource_vector		22'b0000000000000000000000
`define 	vsuxseg3ei32_v_resource_vector		22'b0000000000000000000000
`define 	vsuxseg3ei64_v_resource_vector		22'b0000000000000000000000
`define 	vsuxseg4ei8_v_resource_vector		22'b0000000000000000000000
`define 	vsuxseg4ei16_v_resource_vector		22'b0000000000000000000000
`define 	vsuxseg4ei32_v_resource_vector		22'b0000000000000000000000
`define 	vsuxseg4ei64_v_resource_vector		22'b0000000000000000000000
`define 	vsuxseg5ei8_v_resource_vector		22'b0000000000000000000000
`define 	vsuxseg5ei16_v_resource_vector		22'b0000000000000000000000
`define 	vsuxseg5ei32_v_resource_vector		22'b0000000000000000000000
`define 	vsuxseg5ei64_v_resource_vector		22'b0000000000000000000000
`define 	vsuxseg6ei8_v_resource_vector		22'b0000000000000000000000
`define 	vsuxseg6ei16_v_resource_vector		22'b0000000000000000000000
`define 	vsuxseg6ei32_v_resource_vector		22'b0000000000000000000000
`define 	vsuxseg6ei64_v_resource_vector		22'b0000000000000000000000
`define 	vsuxseg7ei8_v_resource_vector		22'b0000000000000000000000
`define 	vsuxseg7ei16_v_resource_vector		22'b0000000000000000000000
`define 	vsuxseg7ei32_v_resource_vector		22'b0000000000000000000000
`define 	vsuxseg7ei64_v_resource_vector		22'b0000000000000000000000
`define 	vsuxseg8ei8_v_resource_vector		22'b0000000000000000000000
`define 	vsuxseg8ei16_v_resource_vector		22'b0000000000000000000000
`define 	vsuxseg8ei32_v_resource_vector		22'b0000000000000000000000
`define 	vsuxseg8ei64_v_resource_vector		22'b0000000000000000000000
`define 	vsoxseg1ei8_v_resource_vector		22'b0000000000000000000000
`define 	vsoxseg1ei16_v_resource_vector		22'b0000000000000000000000
`define 	vsoxseg1ei32_v_resource_vector		22'b0000000000000000000000
`define 	vsoxseg1ei64_v_resource_vector		22'b0000000000000000000000
`define 	vsoxseg2ei8_v_resource_vector		22'b0000000000000000000000
`define 	vsoxseg2ei16_v_resource_vector		22'b0000000000000000000000
`define 	vsoxseg2ei32_v_resource_vector		22'b0000000000000000000000
`define 	vsoxseg2ei64_v_resource_vector		22'b0000000000000000000000
`define 	vsoxseg3ei8_v_resource_vector		22'b0000000000000000000000
`define 	vsoxseg3ei16_v_resource_vector		22'b0000000000000000000000
`define 	vsoxseg3ei32_v_resource_vector		22'b0000000000000000000000
`define 	vsoxseg3ei64_v_resource_vector		22'b0000000000000000000000
`define 	vsoxseg4ei8_v_resource_vector		22'b0000000000000000000000
`define 	vsoxseg4ei16_v_resource_vector		22'b0000000000000000000000
`define 	vsoxseg4ei32_v_resource_vector		22'b0000000000000000000000
`define 	vsoxseg4ei64_v_resource_vector		22'b0000000000000000000000
`define 	vsoxseg5ei8_v_resource_vector		22'b0000000000000000000000
`define 	vsoxseg5ei16_v_resource_vector		22'b0000000000000000000000
`define 	vsoxseg5ei32_v_resource_vector		22'b0000000000000000000000
`define 	vsoxseg5ei64_v_resource_vector		22'b0000000000000000000000
`define 	vsoxseg6ei8_v_resource_vector		22'b0000000000000000000000
`define 	vsoxseg6ei16_v_resource_vector		22'b0000000000000000000000
`define 	vsoxseg6ei32_v_resource_vector		22'b0000000000000000000000
`define 	vsoxseg6ei64_v_resource_vector		22'b0000000000000000000000
`define 	vsoxseg7ei8_v_resource_vector		22'b0000000000000000000000
`define 	vsoxseg7ei16_v_resource_vector		22'b0000000000000000000000
`define 	vsoxseg7ei32_v_resource_vector		22'b0000000000000000000000
`define 	vsoxseg7ei64_v_resource_vector		22'b0000000000000000000000
`define 	vsoxseg8ei8_v_resource_vector		22'b0000000000000000000000
`define 	vsoxseg8ei16_v_resource_vector		22'b0000000000000000000000
`define 	vsoxseg8ei32_v_resource_vector		22'b0000000000000000000000
`define 	vsoxseg8ei64_v_resource_vector		22'b0000000000000000000000
`define 	vl1re8_v_resource_vector			22'b0000000000000000000000
`define 	vl1re16_v_resource_vector			22'b0000000000000000000000
`define 	vl1re32_v_resource_vector			22'b0000000000000000000000
`define 	vl1re64_v_resource_vector			22'b0000000000000000000000
`define 	vl2re8_v_resource_vector			22'b0000000000000000000000
`define 	vl2re16_v_resource_vector			22'b0000000000000000000000
`define 	vl2re32_v_resource_vector			22'b0000000000000000000000
`define 	vl2re64_v_resource_vector			22'b0000000000000000000000
`define 	vl4re8_v_resource_vector			22'b0000000000000000000000
`define 	vl4re16_v_resource_vector			22'b0000000000000000000000
`define 	vl4re32_v_resource_vector			22'b0000000000000000000000
`define 	vl4re64_v_resource_vector			22'b0000000000000000000000
`define 	vl8re8_v_resource_vector			22'b0000000000000000000000
`define 	vl8re16_v_resource_vector			22'b0000000000000000000000
`define 	vl8re32_v_resource_vector			22'b0000000000000000000000
`define 	vl8re64_v_resource_vector			22'b0000000000000000000000
`define 	vs1r_v_resource_vector				22'b0000000000000000000000
`define 	vs2r_v_resource_vector				22'b0000000000000000000000
`define 	vs4r_v_resource_vector				22'b0000000000000000000000
`define 	vs8r_v_resource_vector				22'b0000000000000000000000

	//register vector
`define 	vle8_v_register_vector				8'b00001100
`define 	vle16_v_register_vector				8'b00001100
`define 	vle32_v_register_vector				8'b00001100
`define 	vle64_v_register_vector				8'b00001100
`define 	vse8_v_register_vector				8'b00010100
`define 	vse16_v_register_vector				8'b00010100
`define 	vse32_v_register_vector				8'b00010100
`define 	vse64_v_register_vector				8'b00010100
`define 	vlm_v_register_vector				8'b00001100
`define 	vsm_v_register_vector				8'b00010100
`define 	vlse8_v_register_vector				8'b00001110
`define 	vlse16_v_register_vector			8'b00001110
`define 	vlse32_v_register_vector			8'b00001110
`define 	vlse64_v_register_vector			8'b00001110
`define 	vsse8_v_register_vector				8'b00010110
`define 	vsse16_v_register_vector			8'b00010110
`define 	vsse32_v_register_vector			8'b00010110
`define 	vsse64_v_register_vector			8'b00010110
`define 	vluxei8_v_register_vector			8'b00101100
`define 	vluxei16_v_register_vector			8'b00101100
`define 	vluxei32_v_register_vector			8'b00101100
`define 	vluxei64_v_register_vector			8'b00101100
`define 	vloxei8_v_register_vector			8'b00101100
`define 	vloxei16_v_register_vector			8'b00101100
`define 	vloxei32_v_register_vector			8'b00101100
`define 	vloxei64_v_register_vector			8'b00101100
`define 	vsuxei8_v_register_vector			8'b00110100
`define 	vsuxei16_v_register_vector			8'b00110100
`define 	vsuxei32_v_register_vector			8'b00110100
`define 	vsuxei64_v_register_vector			8'b00110100
`define 	vsoxei8_v_register_vector			8'b00110100
`define 	vsoxei16_v_register_vector			8'b00110100
`define 	vsoxei32_v_register_vector			8'b00110100
`define 	vsoxei64_v_register_vector			8'b00110100
`define 	vle8ff_v_register_vector			8'b00001100
`define 	vle16ff_v_register_vector			8'b00001100
`define 	vle32ff_v_register_vector			8'b00001100
`define 	vle64ff_v_register_vector			8'b00001100
`define 	vlseg1e8_v_register_vector			8'b00001100
`define 	vlseg1e16_v_register_vector			8'b00001100
`define 	vlseg1e32_v_register_vector			8'b00001100
`define 	vlseg1e64_v_register_vector			8'b00001100
`define 	vlseg2e8_v_register_vector			8'b00001100
`define 	vlseg2e16_v_register_vector			8'b00001100
`define 	vlseg2e32_v_register_vector			8'b00001100
`define 	vlseg2e64_v_register_vector			8'b00001100
`define 	vlseg3e8_v_register_vector			8'b00001100
`define 	vlseg3e16_v_register_vector			8'b00001100
`define 	vlseg3e32_v_register_vector			8'b00001100
`define 	vlseg3e64_v_register_vector			8'b00001100
`define 	vlseg4e8_v_register_vector			8'b00001100
`define 	vlseg4e16_v_register_vector			8'b00001100
`define 	vlseg4e32_v_register_vector			8'b00001100
`define 	vlseg4e64_v_register_vector			8'b00001100
`define 	vlseg5e8_v_register_vector			8'b00001100
`define 	vlseg5e16_v_register_vector			8'b00001100
`define 	vlseg5e32_v_register_vector			8'b00001100
`define 	vlseg5e64_v_register_vector			8'b00001100
`define 	vlseg6e8_v_register_vector			8'b00001100
`define 	vlseg6e16_v_register_vector			8'b00001100
`define 	vlseg6e32_v_register_vector			8'b00001100
`define 	vlseg6e64_v_register_vector			8'b00001100
`define 	vlseg7e8_v_register_vector			8'b00001100
`define 	vlseg7e16_v_register_vector			8'b00001100
`define 	vlseg7e32_v_register_vector			8'b00001100
`define 	vlseg7e64_v_register_vector			8'b00001100
`define 	vlseg8e8_v_register_vector			8'b00001100
`define 	vlseg8e16_v_register_vector			8'b00001100
`define 	vlseg8e32_v_register_vector			8'b00001100
`define 	vlseg8e64_v_register_vector			8'b00001100
`define 	vsseg1e8_v_register_vector			8'b00010100
`define 	vsseg1e16_v_register_vector			8'b00010100
`define 	vsseg1e32_v_register_vector			8'b00010100
`define 	vsseg1e64_v_register_vector			8'b00010100
`define 	vsseg2e8_v_register_vector			8'b00010100
`define 	vsseg2e16_v_register_vector			8'b00010100
`define 	vsseg2e32_v_register_vector			8'b00010100
`define 	vsseg2e64_v_register_vector			8'b00010100
`define 	vsseg3e8_v_register_vector			8'b00010100
`define 	vsseg3e16_v_register_vector			8'b00010100
`define 	vsseg3e32_v_register_vector			8'b00010100
`define 	vsseg3e64_v_register_vector			8'b00010100
`define 	vsseg4e8_v_register_vector			8'b00010100
`define 	vsseg4e16_v_register_vector			8'b00010100
`define 	vsseg4e32_v_register_vector			8'b00010100
`define 	vsseg4e64_v_register_vector			8'b00010100
`define 	vsseg5e8_v_register_vector			8'b00010100
`define 	vsseg5e16_v_register_vector			8'b00010100
`define 	vsseg5e32_v_register_vector			8'b00010100
`define 	vsseg5e64_v_register_vector			8'b00010100
`define 	vsseg6e8_v_register_vector			8'b00010100
`define 	vsseg6e16_v_register_vector			8'b00010100
`define 	vsseg6e32_v_register_vector			8'b00010100
`define 	vsseg6e64_v_register_vector			8'b00010100
`define 	vsseg7e8_v_register_vector			8'b00010100
`define 	vsseg7e16_v_register_vector			8'b00010100
`define 	vsseg7e32_v_register_vector			8'b00010100
`define 	vsseg7e64_v_register_vector			8'b00010100
`define 	vsseg8e8_v_register_vector			8'b00010100
`define 	vsseg8e16_v_register_vector			8'b00010100
`define 	vsseg8e32_v_register_vector			8'b00010100
`define 	vsseg8e64_v_register_vector			8'b00010100
`define 	vlseg1e8ff_v_register_vector		8'b00001100
`define 	vlseg1e16ff_v_register_vector		8'b00001100
`define 	vlseg1e32ff_v_register_vector		8'b00001100
`define 	vlseg1e64ff_v_register_vector		8'b00001100
`define 	vlseg2e8ff_v_register_vector		8'b00001100
`define 	vlseg2e16ff_v_register_vector		8'b00001100
`define 	vlseg2e32ff_v_register_vector		8'b00001100
`define 	vlseg2e64ff_v_register_vector		8'b00001100
`define 	vlseg3e8ff_v_register_vector		8'b00001100
`define 	vlseg3e16ff_v_register_vector		8'b00001100
`define 	vlseg3e32ff_v_register_vector		8'b00001100
`define 	vlseg3e64ff_v_register_vector		8'b00001100
`define 	vlseg4e8ff_v_register_vector		8'b00001100
`define 	vlseg4e16ff_v_register_vector		8'b00001100
`define 	vlseg4e32ff_v_register_vector		8'b00001100
`define 	vlseg4e64ff_v_register_vector		8'b00001100
`define 	vlseg5e8ff_v_register_vector		8'b00001100
`define 	vlseg5e16ff_v_register_vector		8'b00001100
`define 	vlseg5e32ff_v_register_vector		8'b00001100
`define 	vlseg5e64ff_v_register_vector		8'b00001100
`define 	vlseg6e8ff_v_register_vector		8'b00001100
`define 	vlseg6e16ff_v_register_vector		8'b00001100
`define 	vlseg6e32ff_v_register_vector		8'b00001100
`define 	vlseg6e64ff_v_register_vector		8'b00001100
`define 	vlseg7e8ff_v_register_vector		8'b00001100
`define 	vlseg7e16ff_v_register_vector		8'b00001100
`define 	vlseg7e32ff_v_register_vector		8'b00001100
`define 	vlseg7e64ff_v_register_vector		8'b00001100
`define 	vlseg8e8ff_v_register_vector		8'b00001100
`define 	vlseg8e16ff_v_register_vector		8'b00001100
`define 	vlseg8e32ff_v_register_vector		8'b00001100
`define 	vlseg8e64ff_v_register_vector		8'b00001100
`define 	vlsseg1e8_v_register_vector			8'b00001110
`define 	vlsseg1e16_v_register_vector		8'b00001110
`define 	vlsseg1e32_v_register_vector		8'b00001110
`define 	vlsseg1e64_v_register_vector		8'b00001110
`define 	vlsseg2e8_v_register_vector			8'b00001110
`define 	vlsseg2e16_v_register_vector		8'b00001110
`define 	vlsseg2e32_v_register_vector		8'b00001110
`define 	vlsseg2e64_v_register_vector		8'b00001110
`define 	vlsseg3e8_v_register_vector			8'b00001110
`define 	vlsseg3e16_v_register_vector		8'b00001110
`define 	vlsseg3e32_v_register_vector		8'b00001110
`define 	vlsseg3e64_v_register_vector		8'b00001110
`define 	vlsseg4e8_v_register_vector			8'b00001110
`define 	vlsseg4e16_v_register_vector		8'b00001110
`define 	vlsseg4e32_v_register_vector		8'b00001110
`define 	vlsseg4e64_v_register_vector		8'b00001110
`define 	vlsseg5e8_v_register_vector			8'b00001110
`define 	vlsseg5e16_v_register_vector		8'b00001110
`define 	vlsseg5e32_v_register_vector		8'b00001110
`define 	vlsseg5e64_v_register_vector		8'b00001110
`define 	vlsseg6e8_v_register_vector			8'b00001110
`define 	vlsseg6e16_v_register_vector		8'b00001110
`define 	vlsseg6e32_v_register_vector		8'b00001110
`define 	vlsseg6e64_v_register_vector		8'b00001110
`define 	vlsseg7e8_v_register_vector			8'b00001110
`define 	vlsseg7e16_v_register_vector		8'b00001110
`define 	vlsseg7e32_v_register_vector		8'b00001110
`define 	vlsseg7e64_v_register_vector		8'b00001110
`define 	vlsseg8e8_v_register_vector			8'b00001110
`define 	vlsseg8e16_v_register_vector		8'b00001110
`define 	vlsseg8e32_v_register_vector		8'b00001110
`define 	vlsseg8e64_v_register_vector		8'b00001110
`define 	vssseg1e8_v_register_vector			8'b00010110
`define 	vssseg1e16_v_register_vector		8'b00010110
`define 	vssseg1e32_v_register_vector		8'b00010110
`define 	vssseg1e64_v_register_vector		8'b00010110
`define 	vssseg2e8_v_register_vector			8'b00010110
`define 	vssseg2e16_v_register_vector		8'b00010110
`define 	vssseg2e32_v_register_vector		8'b00010110
`define 	vssseg2e64_v_register_vector		8'b00010110
`define 	vssseg3e8_v_register_vector			8'b00010110
`define 	vssseg3e16_v_register_vector		8'b00010110
`define 	vssseg3e32_v_register_vector		8'b00010110
`define 	vssseg3e64_v_register_vector		8'b00010110
`define 	vssseg4e8_v_register_vector			8'b00010110
`define 	vssseg4e16_v_register_vector		8'b00010110
`define 	vssseg4e32_v_register_vector		8'b00010110
`define 	vssseg4e64_v_register_vector		8'b00010110
`define 	vssseg5e8_v_register_vector			8'b00010110
`define 	vssseg5e16_v_register_vector		8'b00010110
`define 	vssseg5e32_v_register_vector		8'b00010110
`define 	vssseg5e64_v_register_vector		8'b00010110
`define 	vssseg6e8_v_register_vector			8'b00010110
`define 	vssseg6e16_v_register_vector		8'b00010110
`define 	vssseg6e32_v_register_vector		8'b00010110
`define 	vssseg6e64_v_register_vector		8'b00010110
`define 	vssseg7e8_v_register_vector			8'b00010110
`define 	vssseg7e16_v_register_vector		8'b00010110
`define 	vssseg7e32_v_register_vector		8'b00010110
`define 	vssseg7e64_v_register_vector		8'b00010110
`define 	vssseg8e8_v_register_vector			8'b00010110
`define 	vssseg8e16_v_register_vector		8'b00010110
`define 	vssseg8e32_v_register_vector		8'b00010110
`define 	vssseg8e64_v_register_vector		8'b00010110
`define 	vluxseg1ei8_v_register_vector		8'b00101100
`define 	vluxseg1ei16_v_register_vector		8'b00101100
`define 	vluxseg1ei32_v_register_vector		8'b00101100
`define 	vluxseg1ei64_v_register_vector		8'b00101100
`define 	vluxseg2ei8_v_register_vector		8'b00101100
`define 	vluxseg2ei16_v_register_vector		8'b00101100
`define 	vluxseg2ei32_v_register_vector		8'b00101100
`define 	vluxseg2ei64_v_register_vector		8'b00101100
`define 	vluxseg3ei8_v_register_vector		8'b00101100
`define 	vluxseg3ei16_v_register_vector		8'b00101100
`define 	vluxseg3ei32_v_register_vector		8'b00101100
`define 	vluxseg3ei64_v_register_vector		8'b00101100
`define 	vluxseg4ei8_v_register_vector		8'b00101100
`define 	vluxseg4ei16_v_register_vector		8'b00101100
`define 	vluxseg4ei32_v_register_vector		8'b00101100
`define 	vluxseg4ei64_v_register_vector		8'b00101100
`define 	vluxseg5ei8_v_register_vector		8'b00101100
`define 	vluxseg5ei16_v_register_vector		8'b00101100
`define 	vluxseg5ei32_v_register_vector		8'b00101100
`define 	vluxseg5ei64_v_register_vector		8'b00101100
`define 	vluxseg6ei8_v_register_vector		8'b00101100
`define 	vluxseg6ei16_v_register_vector		8'b00101100
`define 	vluxseg6ei32_v_register_vector		8'b00101100
`define 	vluxseg6ei64_v_register_vector		8'b00101100
`define 	vluxseg7ei8_v_register_vector		8'b00101100
`define 	vluxseg7ei16_v_register_vector		8'b00101100
`define 	vluxseg7ei32_v_register_vector		8'b00101100
`define 	vluxseg7ei64_v_register_vector		8'b00101100
`define 	vluxseg8ei8_v_register_vector		8'b00101100
`define 	vluxseg8ei16_v_register_vector		8'b00101100
`define 	vluxseg8ei32_v_register_vector		8'b00101100
`define 	vluxseg8ei64_v_register_vector		8'b00101100
`define 	vloxseg1ei8_v_register_vector		8'b00101100
`define 	vloxseg1ei16_v_register_vector		8'b00101100
`define 	vloxseg1ei32_v_register_vector		8'b00101100
`define 	vloxseg1ei64_v_register_vector		8'b00101100
`define 	vloxseg2ei8_v_register_vector		8'b00101100
`define 	vloxseg2ei16_v_register_vector		8'b00101100
`define 	vloxseg2ei32_v_register_vector		8'b00101100
`define 	vloxseg2ei64_v_register_vector		8'b00101100
`define 	vloxseg3ei8_v_register_vector		8'b00101100
`define 	vloxseg3ei16_v_register_vector		8'b00101100
`define 	vloxseg3ei32_v_register_vector		8'b00101100
`define 	vloxseg3ei64_v_register_vector		8'b00101100
`define 	vloxseg4ei8_v_register_vector		8'b00101100
`define 	vloxseg4ei16_v_register_vector		8'b00101100
`define 	vloxseg4ei32_v_register_vector		8'b00101100
`define 	vloxseg4ei64_v_register_vector		8'b00101100
`define 	vloxseg5ei8_v_register_vector		8'b00101100
`define 	vloxseg5ei16_v_register_vector		8'b00101100
`define 	vloxseg5ei32_v_register_vector		8'b00101100
`define 	vloxseg5ei64_v_register_vector		8'b00101100
`define 	vloxseg6ei8_v_register_vector		8'b00101100
`define 	vloxseg6ei16_v_register_vector		8'b00101100
`define 	vloxseg6ei32_v_register_vector		8'b00101100
`define 	vloxseg6ei64_v_register_vector		8'b00101100
`define 	vloxseg7ei8_v_register_vector		8'b00101100
`define 	vloxseg7ei16_v_register_vector		8'b00101100
`define 	vloxseg7ei32_v_register_vector		8'b00101100
`define 	vloxseg7ei64_v_register_vector		8'b00101100
`define 	vloxseg8ei8_v_register_vector		8'b00101100
`define 	vloxseg8ei16_v_register_vector		8'b00101100
`define 	vloxseg8ei32_v_register_vector		8'b00101100
`define 	vloxseg8ei64_v_register_vector		8'b00101100
`define 	vsuxseg1ei8_v_register_vector		8'b00110100
`define 	vsuxseg1ei16_v_register_vector		8'b00110100
`define 	vsuxseg1ei32_v_register_vector		8'b00110100
`define 	vsuxseg1ei64_v_register_vector		8'b00110100
`define 	vsuxseg2ei8_v_register_vector		8'b00110100
`define 	vsuxseg2ei16_v_register_vector		8'b00110100
`define 	vsuxseg2ei32_v_register_vector		8'b00110100
`define 	vsuxseg2ei64_v_register_vector		8'b00110100
`define 	vsuxseg3ei8_v_register_vector		8'b00110100
`define 	vsuxseg3ei16_v_register_vector		8'b00110100
`define 	vsuxseg3ei32_v_register_vector		8'b00110100
`define 	vsuxseg3ei64_v_register_vector		8'b00110100
`define 	vsuxseg4ei8_v_register_vector		8'b00110100
`define 	vsuxseg4ei16_v_register_vector		8'b00110100
`define 	vsuxseg4ei32_v_register_vector		8'b00110100
`define 	vsuxseg4ei64_v_register_vector		8'b00110100
`define 	vsuxseg5ei8_v_register_vector		8'b00110100
`define 	vsuxseg5ei16_v_register_vector		8'b00110100
`define 	vsuxseg5ei32_v_register_vector		8'b00110100
`define 	vsuxseg5ei64_v_register_vector		8'b00110100
`define 	vsuxseg6ei8_v_register_vector		8'b00110100
`define 	vsuxseg6ei16_v_register_vector		8'b00110100
`define 	vsuxseg6ei32_v_register_vector		8'b00110100
`define 	vsuxseg6ei64_v_register_vector		8'b00110100
`define 	vsuxseg7ei8_v_register_vector		8'b00110100
`define 	vsuxseg7ei16_v_register_vector		8'b00110100
`define 	vsuxseg7ei32_v_register_vector		8'b00110100
`define 	vsuxseg7ei64_v_register_vector		8'b00110100
`define 	vsuxseg8ei8_v_register_vector		8'b00110100
`define 	vsuxseg8ei16_v_register_vector		8'b00110100
`define 	vsuxseg8ei32_v_register_vector		8'b00110100
`define 	vsuxseg8ei64_v_register_vector		8'b00110100
`define 	vsoxseg1ei8_v_register_vector		8'b00110100
`define 	vsoxseg1ei16_v_register_vector		8'b00110100
`define 	vsoxseg1ei32_v_register_vector		8'b00110100
`define 	vsoxseg1ei64_v_register_vector		8'b00110100
`define 	vsoxseg2ei8_v_register_vector		8'b00110100
`define 	vsoxseg2ei16_v_register_vector		8'b00110100
`define 	vsoxseg2ei32_v_register_vector		8'b00110100
`define 	vsoxseg2ei64_v_register_vector		8'b00110100
`define 	vsoxseg3ei8_v_register_vector		8'b00110100
`define 	vsoxseg3ei16_v_register_vector		8'b00110100
`define 	vsoxseg3ei32_v_register_vector		8'b00110100
`define 	vsoxseg3ei64_v_register_vector		8'b00110100
`define 	vsoxseg4ei8_v_register_vector		8'b00110100
`define 	vsoxseg4ei16_v_register_vector		8'b00110100
`define 	vsoxseg4ei32_v_register_vector		8'b00110100
`define 	vsoxseg4ei64_v_register_vector		8'b00110100
`define 	vsoxseg5ei8_v_register_vector		8'b00110100
`define 	vsoxseg5ei16_v_register_vector		8'b00110100
`define 	vsoxseg5ei32_v_register_vector		8'b00110100
`define 	vsoxseg5ei64_v_register_vector		8'b00110100
`define 	vsoxseg6ei8_v_register_vector		8'b00110100
`define 	vsoxseg6ei16_v_register_vector		8'b00110100
`define 	vsoxseg6ei32_v_register_vector		8'b00110100
`define 	vsoxseg6ei64_v_register_vector		8'b00110100
`define 	vsoxseg7ei8_v_register_vector		8'b00110100
`define 	vsoxseg7ei16_v_register_vector		8'b00110100
`define 	vsoxseg7ei32_v_register_vector		8'b00110100
`define 	vsoxseg7ei64_v_register_vector		8'b00110100
`define 	vsoxseg8ei8_v_register_vector		8'b00110100
`define 	vsoxseg8ei16_v_register_vector		8'b00110100
`define 	vsoxseg8ei32_v_register_vector		8'b00110100
`define 	vsoxseg8ei64_v_register_vector		8'b00110100
`define 	vl1re8_v_register_vector			8'b00001100
`define 	vl1re16_v_register_vector			8'b00001100
`define 	vl1re32_v_register_vector			8'b00001100
`define 	vl1re64_v_register_vector			8'b00001100
`define 	vl2re8_v_register_vector			8'b00001100
`define 	vl2re16_v_register_vector			8'b00001100
`define 	vl2re32_v_register_vector			8'b00001100
`define 	vl2re64_v_register_vector			8'b00001100
`define 	vl4re8_v_register_vector			8'b00001100
`define 	vl4re16_v_register_vector			8'b00001100
`define 	vl4re32_v_register_vector			8'b00001100
`define 	vl4re64_v_register_vector			8'b00001100
`define 	vl8re8_v_register_vector			8'b00001100
`define 	vl8re16_v_register_vector			8'b00001100
`define 	vl8re32_v_register_vector			8'b00001100
`define 	vl8re64_v_register_vector			8'b00001100
`define 	vs1r_v_register_vector				8'b00010100
`define 	vs2r_v_register_vector				8'b00010100
`define 	vs4r_v_register_vector				8'b00010100
`define 	vs8r_v_register_vector				8'b00010100

	//operation vector
`define 	vle8_v_operation_vector				29'b01011001000100001100000000000
`define 	vle16_v_operation_vector			29'b01011001000100001100000000000
`define 	vle32_v_operation_vector			29'b01011001000100001100000000000
`define 	vle64_v_operation_vector			29'b01011001000100001100000000000
`define 	vse8_v_operation_vector				29'b01011001000100001100000000000
`define 	vse16_v_operation_vector			29'b01011001000100001100000000000
`define 	vse32_v_operation_vector			29'b01011001000100001100000000000
`define 	vse64_v_operation_vector			29'b01011001000100001100000000000
`define 	vlm_v_operation_vector				29'b01010001000100001100000000000
`define 	vsm_v_operation_vector				29'b01010001000100001100000000000
`define 	vlse8_v_operation_vector			29'b01011001000100001100000000000
`define 	vlse16_v_operation_vector			29'b01011001000100001100000000000
`define 	vlse32_v_operation_vector			29'b01011001000100001100000000000
`define 	vlse64_v_operation_vector			29'b01011001000100001100000000000
`define 	vsse8_v_operation_vector			29'b01011001000100001100000000000
`define 	vsse16_v_operation_vector			29'b01011001000100001100000000000
`define 	vsse32_v_operation_vector			29'b01011001000100001100000000000
`define 	vsse64_v_operation_vector			29'b01011001000100001100000000000
`define 	vluxei8_v_operation_vector			29'b01011001000100001100000000000
`define 	vluxei16_v_operation_vector			29'b01011001000100001100000000000
`define 	vluxei32_v_operation_vector			29'b01011001000100001100000000000
`define 	vluxei64_v_operation_vector			29'b01011001000100001100000000000
`define 	vloxei8_v_operation_vector			29'b01011001000100001100000000000
`define 	vloxei16_v_operation_vector			29'b01011001000100001100000000000
`define 	vloxei32_v_operation_vector			29'b01011001000100001100000000000
`define 	vloxei64_v_operation_vector			29'b01011001000100001100000000000
`define 	vsuxei8_v_operation_vector			29'b01011001000100001100000000000
`define 	vsuxei16_v_operation_vector			29'b01011001000100001100000000000
`define 	vsuxei32_v_operation_vector			29'b01011001000100001100000000000
`define 	vsuxei64_v_operation_vector			29'b01011001000100001100000000000
`define 	vsoxei8_v_operation_vector			29'b01011001000100001100000000000
`define 	vsoxei16_v_operation_vector			29'b01011001000100001100000000000
`define 	vsoxei32_v_operation_vector			29'b01011001000100001100000000000
`define 	vsoxei64_v_operation_vector			29'b01011001000100001100000000000
`define 	vle8ff_v_operation_vector			29'b01011001000100001100000000000
`define 	vle16ff_v_operation_vector			29'b01011001000100001100000000000
`define 	vle32ff_v_operation_vector			29'b01011001000100001100000000000
`define 	vle64ff_v_operation_vector			29'b01011001000100001100000000000
`define 	vlseg1e8_v_operation_vector			29'b01011001000100001100000000000
`define 	vlseg1e16_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg1e32_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg1e64_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg2e8_v_operation_vector			29'b01011001000100001100000000000
`define 	vlseg2e16_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg2e32_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg2e64_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg3e8_v_operation_vector			29'b01011001000100001100000000000
`define 	vlseg3e16_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg3e32_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg3e64_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg4e8_v_operation_vector			29'b01011001000100001100000000000
`define 	vlseg4e16_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg4e32_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg4e64_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg5e8_v_operation_vector			29'b01011001000100001100000000000
`define 	vlseg5e16_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg5e32_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg5e64_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg6e8_v_operation_vector			29'b01011001000100001100000000000
`define 	vlseg6e16_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg6e32_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg6e64_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg7e8_v_operation_vector			29'b01011001000100001100000000000
`define 	vlseg7e16_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg7e32_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg7e64_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg8e8_v_operation_vector			29'b01011001000100001100000000000
`define 	vlseg8e16_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg8e32_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg8e64_v_operation_vector		29'b01011001000100001100000000000
`define 	vsseg1e8_v_operation_vector			29'b01011001000100001100000000000
`define 	vsseg1e16_v_operation_vector		29'b01011001000100001100000000000
`define 	vsseg1e32_v_operation_vector		29'b01011001000100001100000000000
`define 	vsseg1e64_v_operation_vector		29'b01011001000100001100000000000
`define 	vsseg2e8_v_operation_vector			29'b01011001000100001100000000000
`define 	vsseg2e16_v_operation_vector		29'b01011001000100001100000000000
`define 	vsseg2e32_v_operation_vector		29'b01011001000100001100000000000
`define 	vsseg2e64_v_operation_vector		29'b01011001000100001100000000000
`define 	vsseg3e8_v_operation_vector			29'b01011001000100001100000000000
`define 	vsseg3e16_v_operation_vector		29'b01011001000100001100000000000
`define 	vsseg3e32_v_operation_vector		29'b01011001000100001100000000000
`define 	vsseg3e64_v_operation_vector		29'b01011001000100001100000000000
`define 	vsseg4e8_v_operation_vector			29'b01011001000100001100000000000
`define 	vsseg4e16_v_operation_vector		29'b01011001000100001100000000000
`define 	vsseg4e32_v_operation_vector		29'b01011001000100001100000000000
`define 	vsseg4e64_v_operation_vector		29'b01011001000100001100000000000
`define 	vsseg5e8_v_operation_vector			29'b01011001000100001100000000000
`define 	vsseg5e16_v_operation_vector		29'b01011001000100001100000000000
`define 	vsseg5e32_v_operation_vector		29'b01011001000100001100000000000
`define 	vsseg5e64_v_operation_vector		29'b01011001000100001100000000000
`define 	vsseg6e8_v_operation_vector			29'b01011001000100001100000000000
`define 	vsseg6e16_v_operation_vector		29'b01011001000100001100000000000
`define 	vsseg6e32_v_operation_vector		29'b01011001000100001100000000000
`define 	vsseg6e64_v_operation_vector		29'b01011001000100001100000000000
`define 	vsseg7e8_v_operation_vector			29'b01011001000100001100000000000
`define 	vsseg7e16_v_operation_vector		29'b01011001000100001100000000000
`define 	vsseg7e32_v_operation_vector		29'b01011001000100001100000000000
`define 	vsseg7e64_v_operation_vector		29'b01011001000100001100000000000
`define 	vsseg8e8_v_operation_vector			29'b01011001000100001100000000000
`define 	vsseg8e16_v_operation_vector		29'b01011001000100001100000000000
`define 	vsseg8e32_v_operation_vector		29'b01011001000100001100000000000
`define 	vsseg8e64_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg1e8ff_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg1e16ff_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg1e32ff_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg1e64ff_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg2e8ff_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg2e16ff_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg2e32ff_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg2e64ff_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg3e8ff_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg3e16ff_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg3e32ff_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg3e64ff_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg4e8ff_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg4e16ff_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg4e32ff_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg4e64ff_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg5e8ff_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg5e16ff_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg5e32ff_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg5e64ff_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg6e8ff_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg6e16ff_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg6e32ff_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg6e64ff_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg7e8ff_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg7e16ff_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg7e32ff_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg7e64ff_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg8e8ff_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg8e16ff_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg8e32ff_v_operation_vector		29'b01011001000100001100000000000
`define 	vlseg8e64ff_v_operation_vector		29'b01011001000100001100000000000
`define 	vlsseg1e8_v_operation_vector		29'b01011001000100001100000000000
`define 	vlsseg1e16_v_operation_vector		29'b01011001000100001100000000000
`define 	vlsseg1e32_v_operation_vector		29'b01011001000100001100000000000
`define 	vlsseg1e64_v_operation_vector		29'b01011001000100001100000000000
`define 	vlsseg2e8_v_operation_vector		29'b01011001000100001100000000000
`define 	vlsseg2e16_v_operation_vector		29'b01011001000100001100000000000
`define 	vlsseg2e32_v_operation_vector		29'b01011001000100001100000000000
`define 	vlsseg2e64_v_operation_vector		29'b01011001000100001100000000000
`define 	vlsseg3e8_v_operation_vector		29'b01011001000100001100000000000
`define 	vlsseg3e16_v_operation_vector		29'b01011001000100001100000000000
`define 	vlsseg3e32_v_operation_vector		29'b01011001000100001100000000000
`define 	vlsseg3e64_v_operation_vector		29'b01011001000100001100000000000
`define 	vlsseg4e8_v_operation_vector		29'b01011001000100001100000000000
`define 	vlsseg4e16_v_operation_vector		29'b01011001000100001100000000000
`define 	vlsseg4e32_v_operation_vector		29'b01011001000100001100000000000
`define 	vlsseg4e64_v_operation_vector		29'b01011001000100001100000000000
`define 	vlsseg5e8_v_operation_vector		29'b01011001000100001100000000000
`define 	vlsseg5e16_v_operation_vector		29'b01011001000100001100000000000
`define 	vlsseg5e32_v_operation_vector		29'b01011001000100001100000000000
`define 	vlsseg5e64_v_operation_vector		29'b01011001000100001100000000000
`define 	vlsseg6e8_v_operation_vector		29'b01011001000100001100000000000
`define 	vlsseg6e16_v_operation_vector		29'b01011001000100001100000000000
`define 	vlsseg6e32_v_operation_vector		29'b01011001000100001100000000000
`define 	vlsseg6e64_v_operation_vector		29'b01011001000100001100000000000
`define 	vlsseg7e8_v_operation_vector		29'b01011001000100001100000000000
`define 	vlsseg7e16_v_operation_vector		29'b01011001000100001100000000000
`define 	vlsseg7e32_v_operation_vector		29'b01011001000100001100000000000
`define 	vlsseg7e64_v_operation_vector		29'b01011001000100001100000000000
`define 	vlsseg8e8_v_operation_vector		29'b01011001000100001100000000000
`define 	vlsseg8e16_v_operation_vector		29'b01011001000100001100000000000
`define 	vlsseg8e32_v_operation_vector		29'b01011001000100001100000000000
`define 	vlsseg8e64_v_operation_vector		29'b01011001000100001100000000000
`define 	vssseg1e8_v_operation_vector		29'b01011001000100001100000000000
`define 	vssseg1e16_v_operation_vector		29'b01011001000100001100000000000
`define 	vssseg1e32_v_operation_vector		29'b01011001000100001100000000000
`define 	vssseg1e64_v_operation_vector		29'b01011001000100001100000000000
`define 	vssseg2e8_v_operation_vector		29'b01011001000100001100000000000
`define 	vssseg2e16_v_operation_vector		29'b01011001000100001100000000000
`define 	vssseg2e32_v_operation_vector		29'b01011001000100001100000000000
`define 	vssseg2e64_v_operation_vector		29'b01011001000100001100000000000
`define 	vssseg3e8_v_operation_vector		29'b01011001000100001100000000000
`define 	vssseg3e16_v_operation_vector		29'b01011001000100001100000000000
`define 	vssseg3e32_v_operation_vector		29'b01011001000100001100000000000
`define 	vssseg3e64_v_operation_vector		29'b01011001000100001100000000000
`define 	vssseg4e8_v_operation_vector		29'b01011001000100001100000000000
`define 	vssseg4e16_v_operation_vector		29'b01011001000100001100000000000
`define 	vssseg4e32_v_operation_vector		29'b01011001000100001100000000000
`define 	vssseg4e64_v_operation_vector		29'b01011001000100001100000000000
`define 	vssseg5e8_v_operation_vector		29'b01011001000100001100000000000
`define 	vssseg5e16_v_operation_vector		29'b01011001000100001100000000000
`define 	vssseg5e32_v_operation_vector		29'b01011001000100001100000000000
`define 	vssseg5e64_v_operation_vector		29'b01011001000100001100000000000
`define 	vssseg6e8_v_operation_vector		29'b01011001000100001100000000000
`define 	vssseg6e16_v_operation_vector		29'b01011001000100001100000000000
`define 	vssseg6e32_v_operation_vector		29'b01011001000100001100000000000
`define 	vssseg6e64_v_operation_vector		29'b01011001000100001100000000000
`define 	vssseg7e8_v_operation_vector		29'b01011001000100001100000000000
`define 	vssseg7e16_v_operation_vector		29'b01011001000100001100000000000
`define 	vssseg7e32_v_operation_vector		29'b01011001000100001100000000000
`define 	vssseg7e64_v_operation_vector		29'b01011001000100001100000000000
`define 	vssseg8e8_v_operation_vector		29'b01011001000100001100000000000
`define 	vssseg8e16_v_operation_vector		29'b01011001000100001100000000000
`define 	vssseg8e32_v_operation_vector		29'b01011001000100001100000000000
`define 	vssseg8e64_v_operation_vector		29'b01011001000100001100000000000
`define 	vluxseg1ei8_v_operation_vector		29'b01011001000100001100000000000
`define 	vluxseg1ei16_v_operation_vector		29'b01011001000100001100000000000
`define 	vluxseg1ei32_v_operation_vector		29'b01011001000100001100000000000
`define 	vluxseg1ei64_v_operation_vector		29'b01011001000100001100000000000
`define 	vluxseg2ei8_v_operation_vector		29'b01011001000100001100000000000
`define 	vluxseg2ei16_v_operation_vector		29'b01011001000100001100000000000
`define 	vluxseg2ei32_v_operation_vector		29'b01011001000100001100000000000
`define 	vluxseg2ei64_v_operation_vector		29'b01011001000100001100000000000
`define 	vluxseg3ei8_v_operation_vector		29'b01011001000100001100000000000
`define 	vluxseg3ei16_v_operation_vector		29'b01011001000100001100000000000
`define 	vluxseg3ei32_v_operation_vector		29'b01011001000100001100000000000
`define 	vluxseg3ei64_v_operation_vector		29'b01011001000100001100000000000
`define 	vluxseg4ei8_v_operation_vector		29'b01011001000100001100000000000
`define 	vluxseg4ei16_v_operation_vector		29'b01011001000100001100000000000
`define 	vluxseg4ei32_v_operation_vector		29'b01011001000100001100000000000
`define 	vluxseg4ei64_v_operation_vector		29'b01011001000100001100000000000
`define 	vluxseg5ei8_v_operation_vector		29'b01011001000100001100000000000
`define 	vluxseg5ei16_v_operation_vector		29'b01011001000100001100000000000
`define 	vluxseg5ei32_v_operation_vector		29'b01011001000100001100000000000
`define 	vluxseg5ei64_v_operation_vector		29'b01011001000100001100000000000
`define 	vluxseg6ei8_v_operation_vector		29'b01011001000100001100000000000
`define 	vluxseg6ei16_v_operation_vector		29'b01011001000100001100000000000
`define 	vluxseg6ei32_v_operation_vector		29'b01011001000100001100000000000
`define 	vluxseg6ei64_v_operation_vector		29'b01011001000100001100000000000
`define 	vluxseg7ei8_v_operation_vector		29'b01011001000100001100000000000
`define 	vluxseg7ei16_v_operation_vector		29'b01011001000100001100000000000
`define 	vluxseg7ei32_v_operation_vector		29'b01011001000100001100000000000
`define 	vluxseg7ei64_v_operation_vector		29'b01011001000100001100000000000
`define 	vluxseg8ei8_v_operation_vector		29'b01011001000100001100000000000
`define 	vluxseg8ei16_v_operation_vector		29'b01011001000100001100000000000
`define 	vluxseg8ei32_v_operation_vector		29'b01011001000100001100000000000
`define 	vluxseg8ei64_v_operation_vector		29'b01011001000100001100000000000
`define 	vloxseg1ei8_v_operation_vector		29'b01011001000100001100000000000
`define 	vloxseg1ei16_v_operation_vector		29'b01011001000100001100000000000
`define 	vloxseg1ei32_v_operation_vector		29'b01011001000100001100000000000
`define 	vloxseg1ei64_v_operation_vector		29'b01011001000100001100000000000
`define 	vloxseg2ei8_v_operation_vector		29'b01011001000100001100000000000
`define 	vloxseg2ei16_v_operation_vector		29'b01011001000100001100000000000
`define 	vloxseg2ei32_v_operation_vector		29'b01011001000100001100000000000
`define 	vloxseg2ei64_v_operation_vector		29'b01011001000100001100000000000
`define 	vloxseg3ei8_v_operation_vector		29'b01011001000100001100000000000
`define 	vloxseg3ei16_v_operation_vector		29'b01011001000100001100000000000
`define 	vloxseg3ei32_v_operation_vector		29'b01011001000100001100000000000
`define 	vloxseg3ei64_v_operation_vector		29'b01011001000100001100000000000
`define 	vloxseg4ei8_v_operation_vector		29'b01011001000100001100000000000
`define 	vloxseg4ei16_v_operation_vector		29'b01011001000100001100000000000
`define 	vloxseg4ei32_v_operation_vector		29'b01011001000100001100000000000
`define 	vloxseg4ei64_v_operation_vector		29'b01011001000100001100000000000
`define 	vloxseg5ei8_v_operation_vector		29'b01011001000100001100000000000
`define 	vloxseg5ei16_v_operation_vector		29'b01011001000100001100000000000
`define 	vloxseg5ei32_v_operation_vector		29'b01011001000100001100000000000
`define 	vloxseg5ei64_v_operation_vector		29'b01011001000100001100000000000
`define 	vloxseg6ei8_v_operation_vector		29'b01011001000100001100000000000
`define 	vloxseg6ei16_v_operation_vector		29'b01011001000100001100000000000
`define 	vloxseg6ei32_v_operation_vector		29'b01011001000100001100000000000
`define 	vloxseg6ei64_v_operation_vector		29'b01011001000100001100000000000
`define 	vloxseg7ei8_v_operation_vector		29'b01011001000100001100000000000
`define 	vloxseg7ei16_v_operation_vector		29'b01011001000100001100000000000
`define 	vloxseg7ei32_v_operation_vector		29'b01011001000100001100000000000
`define 	vloxseg7ei64_v_operation_vector		29'b01011001000100001100000000000
`define 	vloxseg8ei8_v_operation_vector		29'b01011001000100001100000000000
`define 	vloxseg8ei16_v_operation_vector		29'b01011001000100001100000000000
`define 	vloxseg8ei32_v_operation_vector		29'b01011001000100001100000000000
`define 	vloxseg8ei64_v_operation_vector		29'b01011001000100001100000000000
`define 	vsuxseg1ei8_v_operation_vector		29'b01011001000100001100000000000
`define 	vsuxseg1ei16_v_operation_vector		29'b01011001000100001100000000000
`define 	vsuxseg1ei32_v_operation_vector		29'b01011001000100001100000000000
`define 	vsuxseg1ei64_v_operation_vector		29'b01011001000100001100000000000
`define 	vsuxseg2ei8_v_operation_vector		29'b01011001000100001100000000000
`define 	vsuxseg2ei16_v_operation_vector		29'b01011001000100001100000000000
`define 	vsuxseg2ei32_v_operation_vector		29'b01011001000100001100000000000
`define 	vsuxseg2ei64_v_operation_vector		29'b01011001000100001100000000000
`define 	vsuxseg3ei8_v_operation_vector		29'b01011001000100001100000000000
`define 	vsuxseg3ei16_v_operation_vector		29'b01011001000100001100000000000
`define 	vsuxseg3ei32_v_operation_vector		29'b01011001000100001100000000000
`define 	vsuxseg3ei64_v_operation_vector		29'b01011001000100001100000000000
`define 	vsuxseg4ei8_v_operation_vector		29'b01011001000100001100000000000
`define 	vsuxseg4ei16_v_operation_vector		29'b01011001000100001100000000000
`define 	vsuxseg4ei32_v_operation_vector		29'b01011001000100001100000000000
`define 	vsuxseg4ei64_v_operation_vector		29'b01011001000100001100000000000
`define 	vsuxseg5ei8_v_operation_vector		29'b01011001000100001100000000000
`define 	vsuxseg5ei16_v_operation_vector		29'b01011001000100001100000000000
`define 	vsuxseg5ei32_v_operation_vector		29'b01011001000100001100000000000
`define 	vsuxseg5ei64_v_operation_vector		29'b01011001000100001100000000000
`define 	vsuxseg6ei8_v_operation_vector		29'b01011001000100001100000000000
`define 	vsuxseg6ei16_v_operation_vector		29'b01011001000100001100000000000
`define 	vsuxseg6ei32_v_operation_vector		29'b01011001000100001100000000000
`define 	vsuxseg6ei64_v_operation_vector		29'b01011001000100001100000000000
`define 	vsuxseg7ei8_v_operation_vector		29'b01011001000100001100000000000
`define 	vsuxseg7ei16_v_operation_vector		29'b01011001000100001100000000000
`define 	vsuxseg7ei32_v_operation_vector		29'b01011001000100001100000000000
`define 	vsuxseg7ei64_v_operation_vector		29'b01011001000100001100000000000
`define 	vsuxseg8ei8_v_operation_vector		29'b01011001000100001100000000000
`define 	vsuxseg8ei16_v_operation_vector		29'b01011001000100001100000000000
`define 	vsuxseg8ei32_v_operation_vector		29'b01011001000100001100000000000
`define 	vsuxseg8ei64_v_operation_vector		29'b01011001000100001100000000000
`define 	vsoxseg1ei8_v_operation_vector		29'b01011001000100001100000000000
`define 	vsoxseg1ei16_v_operation_vector		29'b01011001000100001100000000000
`define 	vsoxseg1ei32_v_operation_vector		29'b01011001000100001100000000000
`define 	vsoxseg1ei64_v_operation_vector		29'b01011001000100001100000000000
`define 	vsoxseg2ei8_v_operation_vector		29'b01011001000100001100000000000
`define 	vsoxseg2ei16_v_operation_vector		29'b01011001000100001100000000000
`define 	vsoxseg2ei32_v_operation_vector		29'b01011001000100001100000000000
`define 	vsoxseg2ei64_v_operation_vector		29'b01011001000100001100000000000
`define 	vsoxseg3ei8_v_operation_vector		29'b01011001000100001100000000000
`define 	vsoxseg3ei16_v_operation_vector		29'b01011001000100001100000000000
`define 	vsoxseg3ei32_v_operation_vector		29'b01011001000100001100000000000
`define 	vsoxseg3ei64_v_operation_vector		29'b01011001000100001100000000000
`define 	vsoxseg4ei8_v_operation_vector		29'b01011001000100001100000000000
`define 	vsoxseg4ei16_v_operation_vector		29'b01011001000100001100000000000
`define 	vsoxseg4ei32_v_operation_vector		29'b01011001000100001100000000000
`define 	vsoxseg4ei64_v_operation_vector		29'b01011001000100001100000000000
`define 	vsoxseg5ei8_v_operation_vector		29'b01011001000100001100000000000
`define 	vsoxseg5ei16_v_operation_vector		29'b01011001000100001100000000000
`define 	vsoxseg5ei32_v_operation_vector		29'b01011001000100001100000000000
`define 	vsoxseg5ei64_v_operation_vector		29'b01011001000100001100000000000
`define 	vsoxseg6ei8_v_operation_vector		29'b01011001000100001100000000000
`define 	vsoxseg6ei16_v_operation_vector		29'b01011001000100001100000000000
`define 	vsoxseg6ei32_v_operation_vector		29'b01011001000100001100000000000
`define 	vsoxseg6ei64_v_operation_vector		29'b01011001000100001100000000000
`define 	vsoxseg7ei8_v_operation_vector		29'b01011001000100001100000000000
`define 	vsoxseg7ei16_v_operation_vector		29'b01011001000100001100000000000
`define 	vsoxseg7ei32_v_operation_vector		29'b01011001000100001100000000000
`define 	vsoxseg7ei64_v_operation_vector		29'b01011001000100001100000000000
`define 	vsoxseg8ei8_v_operation_vector		29'b01011001000100001100000000000
`define 	vsoxseg8ei16_v_operation_vector		29'b01011001000100001100000000000
`define 	vsoxseg8ei32_v_operation_vector		29'b01011001000100001100000000000
`define 	vsoxseg8ei64_v_operation_vector		29'b01011001000100001100000000000
`define 	vl1re8_v_operation_vector			29'b01011001000100001100000000000
`define 	vl1re16_v_operation_vector			29'b01011001000100001100000000000
`define 	vl1re32_v_operation_vector			29'b01011001000100001100000000000
`define 	vl1re64_v_operation_vector			29'b01011001000100001100000000000
`define 	vl2re8_v_operation_vector			29'b01011001000100001100000000000
`define 	vl2re16_v_operation_vector			29'b01011001000100001100000000000
`define 	vl2re32_v_operation_vector			29'b01011001000100001100000000000
`define 	vl2re64_v_operation_vector			29'b01011001000100001100000000000
`define 	vl4re8_v_operation_vector			29'b01011001000100001100000000000
`define 	vl4re16_v_operation_vector			29'b01011001000100001100000000000
`define 	vl4re32_v_operation_vector			29'b01011001000100001100000000000
`define 	vl4re64_v_operation_vector			29'b01011001000100001100000000000
`define 	vl8re8_v_operation_vector			29'b01011001000100001100000000000
`define 	vl8re16_v_operation_vector			29'b01011001000100001100000000000
`define 	vl8re32_v_operation_vector			29'b01011001000100001100000000000
`define 	vl8re64_v_operation_vector			29'b01011001000100001100000000000
`define 	vs1r_v_operation_vector				29'b01011001000100001100000000000
`define 	vs2r_v_operation_vector				29'b01011001000100001100000000000
`define 	vs4r_v_operation_vector				29'b01011001000100001100000000000
`define 	vs8r_v_operation_vector				29'b01011001000100001100000000000